
module RR_arbiter ( clk, rst, req, gnt );
  input [15:0] req;
  output [15:0] gnt;
  input clk, rst;
  wire   \req_vec_rr[0][3] , \req_vec_rr[0][2] , \req_vec_rr[0][1] ,
         \req_vec_rr[0][0] , \req_vec_rr[1][3] , \req_vec_rr[1][2] ,
         \req_vec_rr[1][1] , \req_vec_rr[1][0] , \req_vec_rr[2][2] ,
         \req_vec_rr[2][1] , \req_vec_rr[2][0] , \req_vec_rr[3][3] ,
         \req_vec_rr[3][2] , \req_vec_rr[3][1] , \req_vec_rr[3][0] ,
         \req_vec_rr[4][3] , \req_vec_rr[4][2] , \req_vec_rr[4][1] ,
         \req_vec_rr[4][0] , \req_vec_rr[5][3] , \req_vec_rr[5][2] ,
         \req_vec_rr[5][1] , \req_vec_rr[5][0] , \req_vec_rr[6][3] ,
         \req_vec_rr[6][2] , \req_vec_rr[6][1] , \req_vec_rr[6][0] ,
         \req_vec_rr[7][3] , \req_vec_rr[7][2] , \req_vec_rr[7][1] ,
         \req_vec_rr[7][0] , \req_vec_rr[8][3] , \req_vec_rr[8][2] ,
         \req_vec_rr[8][1] , \req_vec_rr[8][0] , \req_vec_rr[9][3] ,
         \req_vec_rr[9][2] , \req_vec_rr[9][1] , \req_vec_rr[9][0] ,
         \req_vec_rr[10][3] , \req_vec_rr[10][2] , \req_vec_rr[10][1] ,
         \req_vec_rr[10][0] , \req_vec_rr[11][3] , \req_vec_rr[11][2] ,
         \req_vec_rr[11][1] , \req_vec_rr[11][0] , \req_vec_rr[12][3] ,
         \req_vec_rr[12][2] , \req_vec_rr[12][1] , \req_vec_rr[12][0] ,
         \req_vec_rr[13][3] , \req_vec_rr[13][2] , \req_vec_rr[13][1] ,
         \req_vec_rr[13][0] , \req_vec_rr[14][2] , \req_vec_rr[14][1] ,
         \req_vec_rr[14][0] , \req_vec_rr[15][3] , \req_vec_rr[15][2] ,
         \req_vec_rr[15][1] , \req_vec_rr[15][0] , \req_vec_rr_d[0][3] ,
         \req_vec_rr_d[0][2] , \req_vec_rr_d[0][1] , \req_vec_rr_d[0][0] ,
         \req_vec_rr_d[1][3] , \req_vec_rr_d[1][2] , \req_vec_rr_d[1][1] ,
         \req_vec_rr_d[2][2] , \req_vec_rr_d[2][1] , \req_vec_rr_d[2][0] ,
         \req_vec_rr_d[3][3] , \req_vec_rr_d[3][2] , \req_vec_rr_d[4][3] ,
         \req_vec_rr_d[4][2] , \req_vec_rr_d[4][1] , \req_vec_rr_d[4][0] ,
         \req_vec_rr_d[5][3] , \req_vec_rr_d[5][2] , \req_vec_rr_d[5][1] ,
         \req_vec_rr_d[6][3] , \req_vec_rr_d[6][2] , \req_vec_rr_d[6][1] ,
         \req_vec_rr_d[6][0] , \req_vec_rr_d[7][3] , \req_vec_rr_d[8][3] ,
         \req_vec_rr_d[8][2] , \req_vec_rr_d[8][1] , \req_vec_rr_d[8][0] ,
         \req_vec_rr_d[9][3] , \req_vec_rr_d[9][2] , \req_vec_rr_d[9][1] ,
         \req_vec_rr_d[10][3] , \req_vec_rr_d[10][2] , \req_vec_rr_d[10][1] ,
         \req_vec_rr_d[10][0] , \req_vec_rr_d[11][3] , \req_vec_rr_d[11][2] ,
         \req_vec_rr_d[12][3] , \req_vec_rr_d[12][2] , \req_vec_rr_d[12][1] ,
         \req_vec_rr_d[12][0] , \req_vec_rr_d[13][3] , \req_vec_rr_d[13][2] ,
         \req_vec_rr_d[13][1] , \req_vec_rr_d[14][3] , \req_vec_rr_d[14][2] ,
         \req_vec_rr_d[14][1] , \req_vec_rr_d[14][0] , \req_vec_rr_d[15][3] ,
         \req_vec_rr_d[15][2] , \req_vec_rr_d[15][1] , \req_vec_rr_d[15][0] ,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2403, n2404, n2405, n2406,
         n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416,
         n2417, n2418, n2419, n2420, n2421;
  wire   [15:0] gnt_nxt;

  CFD4QXL \req_vec_rr_reg[15][2]  ( .D(\req_vec_rr_d[15][2] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[15][2] ) );
  CFD4QXL \req_vec_rr_reg[14][2]  ( .D(\req_vec_rr_d[14][2] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[14][2] ) );
  CFD2QX1 \req_vec_rr_reg[9][2]  ( .D(\req_vec_rr_d[9][2] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[9][2] ) );
  CFD2QX1 \req_vec_rr_reg[6][3]  ( .D(\req_vec_rr_d[6][3] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[6][3] ) );
  CFD2QX1 \req_vec_rr_reg[4][3]  ( .D(\req_vec_rr_d[4][3] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[4][3] ) );
  CFD2QX1 \req_vec_rr_reg[3][3]  ( .D(\req_vec_rr_d[3][3] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[3][3] ) );
  CFD2QX1 \req_vec_rr_reg[1][3]  ( .D(\req_vec_rr_d[1][3] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[1][3] ) );
  CFD4QX4 \req_vec_rr_reg[3][1]  ( .D(n2410), .CP(clk), .SD(n2412), .Q(
        \req_vec_rr[3][1] ) );
  CFD2QX4 \req_vec_rr_reg[8][1]  ( .D(\req_vec_rr_d[8][1] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[8][1] ) );
  CFD2QX2 \req_vec_rr_reg[1][2]  ( .D(\req_vec_rr_d[1][2] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[1][2] ) );
  CFD2QX4 \req_vec_rr_reg[4][1]  ( .D(\req_vec_rr_d[4][1] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[4][1] ) );
  CFD2QXL \gnt_d_reg[11]  ( .D(gnt_nxt[11]), .CP(clk), .CD(n2412), .Q(gnt[11])
         );
  CFD2QXL \gnt_d_reg[15]  ( .D(gnt_nxt[15]), .CP(clk), .CD(n2412), .Q(gnt[15])
         );
  CFD2QXL \gnt_d_reg[2]  ( .D(gnt_nxt[2]), .CP(clk), .CD(n2412), .Q(gnt[2]) );
  CFD2QXL \gnt_d_reg[6]  ( .D(gnt_nxt[6]), .CP(clk), .CD(n2412), .Q(gnt[6]) );
  CFD2QXL \gnt_d_reg[3]  ( .D(gnt_nxt[3]), .CP(clk), .CD(n2412), .Q(gnt[3]) );
  CFD2QXL \gnt_d_reg[5]  ( .D(gnt_nxt[5]), .CP(clk), .CD(n2412), .Q(gnt[5]) );
  CFD2QXL \gnt_d_reg[7]  ( .D(gnt_nxt[7]), .CP(clk), .CD(n2412), .Q(gnt[7]) );
  CFD2QXL \gnt_d_reg[8]  ( .D(gnt_nxt[8]), .CP(clk), .CD(n2412), .Q(gnt[8]) );
  CFD2QXL \gnt_d_reg[10]  ( .D(gnt_nxt[10]), .CP(clk), .CD(n2412), .Q(gnt[10])
         );
  CFD2QXL \gnt_d_reg[14]  ( .D(gnt_nxt[14]), .CP(clk), .CD(n2412), .Q(gnt[14])
         );
  CFD2QXL \gnt_d_reg[9]  ( .D(gnt_nxt[9]), .CP(clk), .CD(n2412), .Q(gnt[9]) );
  CFD2QXL \gnt_d_reg[13]  ( .D(gnt_nxt[13]), .CP(clk), .CD(n2412), .Q(gnt[13])
         );
  CFD4QX1 \req_vec_rr_reg[15][3]  ( .D(\req_vec_rr_d[15][3] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[15][3] ) );
  CFD4QX1 \req_vec_rr_reg[11][3]  ( .D(\req_vec_rr_d[11][3] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[11][3] ) );
  CFD4QX1 \req_vec_rr_reg[14][1]  ( .D(\req_vec_rr_d[14][1] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[14][1] ) );
  CFD4QX1 \req_vec_rr_reg[13][2]  ( .D(\req_vec_rr_d[13][2] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[13][2] ) );
  CFD4QX1 \req_vec_rr_reg[11][1]  ( .D(n2411), .CP(clk), .SD(n2412), .Q(
        \req_vec_rr[11][1] ) );
  CFD4QX1 \req_vec_rr_reg[10][1]  ( .D(\req_vec_rr_d[10][1] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[10][1] ) );
  CFD4QX1 \req_vec_rr_reg[12][2]  ( .D(\req_vec_rr_d[12][2] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[12][2] ) );
  CFD4QX2 \req_vec_rr_reg[2][1]  ( .D(\req_vec_rr_d[2][1] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[2][1] ) );
  CFD4QX2 \req_vec_rr_reg[7][1]  ( .D(n2409), .CP(clk), .SD(n2412), .Q(
        \req_vec_rr[7][1] ) );
  CFD4QX1 \req_vec_rr_reg[4][2]  ( .D(\req_vec_rr_d[4][2] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[4][2] ) );
  CFD4QX2 \req_vec_rr_reg[15][0]  ( .D(\req_vec_rr_d[15][0] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[15][0] ) );
  CFD2QX1 \req_vec_rr_reg[0][2]  ( .D(\req_vec_rr_d[0][2] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[0][2] ) );
  CFD2QXL \req_vec_rr_reg[0][3]  ( .D(\req_vec_rr_d[0][3] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[0][3] ) );
  CFD4QX4 \req_vec_rr_reg[6][2]  ( .D(\req_vec_rr_d[6][2] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[6][2] ) );
  CFD2QX2 \req_vec_rr_reg[14][0]  ( .D(\req_vec_rr_d[14][0] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[14][0] ) );
  CFD2QX4 \req_vec_rr_reg[12][0]  ( .D(\req_vec_rr_d[12][0] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[12][0] ) );
  CFD2QX2 \req_vec_rr_reg[7][3]  ( .D(\req_vec_rr_d[7][3] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[7][3] ) );
  CFD2QX2 \req_vec_rr_reg[0][0]  ( .D(\req_vec_rr_d[0][0] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[0][0] ) );
  CFD2QX4 \req_vec_rr_reg[1][1]  ( .D(\req_vec_rr_d[1][1] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[1][1] ) );
  CFD2QX2 \req_vec_rr_reg[5][1]  ( .D(\req_vec_rr_d[5][1] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[5][1] ) );
  CFD2QX2 \req_vec_rr_reg[11][2]  ( .D(\req_vec_rr_d[11][2] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[11][2] ) );
  CFD2QX2 \req_vec_rr_reg[3][2]  ( .D(\req_vec_rr_d[3][2] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[3][2] ) );
  CFD2QX2 \req_vec_rr_reg[12][1]  ( .D(\req_vec_rr_d[12][1] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[12][1] ) );
  CFD4QX2 \req_vec_rr_reg[13][3]  ( .D(\req_vec_rr_d[13][3] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[13][3] ) );
  CFD4QX2 \req_vec_rr_reg[5][2]  ( .D(\req_vec_rr_d[5][2] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[5][2] ) );
  CFD4X1 \req_vec_rr_reg[7][2]  ( .D(n2406), .CP(clk), .SD(n2412), .Q(
        \req_vec_rr[7][2] ), .QN(n2415) );
  CFD4X1 \req_vec_rr_reg[8][3]  ( .D(\req_vec_rr_d[8][3] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[8][3] ), .QN(n2414) );
  CFD4X1 \req_vec_rr_reg[12][3]  ( .D(\req_vec_rr_d[12][3] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[12][3] ), .QN(n2413) );
  CFD4X1 \req_vec_rr_reg[10][3]  ( .D(\req_vec_rr_d[10][3] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[10][3] ), .QN(n2416) );
  CFD4QX2 \req_vec_rr_reg[6][1]  ( .D(\req_vec_rr_d[6][1] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[6][1] ) );
  CFD2QX4 \req_vec_rr_reg[13][1]  ( .D(\req_vec_rr_d[13][1] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[13][1] ) );
  CFD4X1 \req_vec_rr_reg[14][3]  ( .D(\req_vec_rr_d[14][3] ), .CP(clk), .SD(
        n2412), .Q(n2403), .QN(n2404) );
  CFD2XL \gnt_d_reg[12]  ( .D(gnt_nxt[12]), .CP(clk), .CD(n2412), .Q(gnt[12])
         );
  CFD2XL \gnt_d_reg[0]  ( .D(gnt_nxt[0]), .CP(clk), .CD(n2412), .Q(gnt[0]) );
  CFD2XL \gnt_d_reg[4]  ( .D(gnt_nxt[4]), .CP(clk), .CD(n2412), .Q(gnt[4]) );
  CFD2XL \gnt_d_reg[1]  ( .D(gnt_nxt[1]), .CP(clk), .CD(n2412), .Q(gnt[1]) );
  CFD3QX2 \req_vec_rr_reg[11][0]  ( .D(n2407), .CP(clk), .CD(1'b1), .SD(n2412), 
        .Q(\req_vec_rr[11][0] ) );
  CFD3QX2 \req_vec_rr_reg[15][1]  ( .D(\req_vec_rr_d[15][1] ), .CP(clk), .CD(
        1'b1), .SD(n2412), .Q(\req_vec_rr[15][1] ) );
  CFD2QX4 \req_vec_rr_reg[8][2]  ( .D(\req_vec_rr_d[8][2] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[8][2] ) );
  CFD2QX2 \req_vec_rr_reg[5][3]  ( .D(\req_vec_rr_d[5][3] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[5][3] ) );
  CFD2QX4 \req_vec_rr_reg[10][0]  ( .D(\req_vec_rr_d[10][0] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[10][0] ) );
  CFD4QX4 \req_vec_rr_reg[1][0]  ( .D(n2405), .CP(clk), .SD(n2412), .Q(
        \req_vec_rr[1][0] ) );
  CFD2QX4 \req_vec_rr_reg[2][0]  ( .D(\req_vec_rr_d[2][0] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[2][0] ) );
  CFD2QX4 \req_vec_rr_reg[4][0]  ( .D(\req_vec_rr_d[4][0] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[4][0] ) );
  CFD2QX4 \req_vec_rr_reg[8][0]  ( .D(\req_vec_rr_d[8][0] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[8][0] ) );
  CFD2X1 \req_vec_rr_reg[2][3]  ( .D(n2417), .CP(clk), .CD(n2412), .Q(n933), 
        .QN(n932) );
  CFD4QX1 \req_vec_rr_reg[5][0]  ( .D(n2420), .CP(clk), .SD(n2412), .Q(
        \req_vec_rr[5][0] ) );
  CFD4QX1 \req_vec_rr_reg[9][0]  ( .D(n2408), .CP(clk), .SD(n2412), .Q(
        \req_vec_rr[9][0] ) );
  CFD4QX1 \req_vec_rr_reg[3][0]  ( .D(n2421), .CP(clk), .SD(n2412), .Q(
        \req_vec_rr[3][0] ) );
  CFD4QX2 \req_vec_rr_reg[13][0]  ( .D(n2418), .CP(clk), .SD(n2412), .Q(
        \req_vec_rr[13][0] ) );
  CFD4QX2 \req_vec_rr_reg[7][0]  ( .D(n2419), .CP(clk), .SD(n2412), .Q(
        \req_vec_rr[7][0] ) );
  CFD2QX2 \req_vec_rr_reg[6][0]  ( .D(\req_vec_rr_d[6][0] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[6][0] ) );
  CFD2QX2 \req_vec_rr_reg[9][1]  ( .D(\req_vec_rr_d[9][1] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[9][1] ) );
  CFD4QX2 \req_vec_rr_reg[9][3]  ( .D(\req_vec_rr_d[9][3] ), .CP(clk), .SD(
        n2412), .Q(\req_vec_rr[9][3] ) );
  CFD2QX4 \req_vec_rr_reg[2][2]  ( .D(\req_vec_rr_d[2][2] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[2][2] ) );
  CFD2QX4 \req_vec_rr_reg[10][2]  ( .D(\req_vec_rr_d[10][2] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[10][2] ) );
  CFD2QX4 \req_vec_rr_reg[0][1]  ( .D(\req_vec_rr_d[0][1] ), .CP(clk), .CD(
        n2412), .Q(\req_vec_rr[0][1] ) );
  CND2X4 U910 ( .A(n1309), .B(n1308), .Z(n1460) );
  CNR2X4 U911 ( .A(n2273), .B(n2300), .Z(n1742) );
  CND2X2 U912 ( .A(n909), .B(n907), .Z(n1980) );
  CIVX2 U913 ( .A(n908), .Z(n907) );
  CND2X2 U914 ( .A(n914), .B(n1905), .Z(n908) );
  CIVX1 U915 ( .A(n2291), .Z(n909) );
  CNR2IX2 U916 ( .B(n1905), .A(n2291), .Z(n916) );
  CND2X2 U917 ( .A(n916), .B(n910), .Z(n1472) );
  CIVX2 U918 ( .A(n911), .Z(n910) );
  CND2X2 U919 ( .A(n1972), .B(n1794), .Z(n911) );
  CND2X2 U920 ( .A(n916), .B(n912), .Z(n1931) );
  CIVX2 U921 ( .A(n913), .Z(n912) );
  CND2X2 U922 ( .A(n2293), .B(n2018), .Z(n913) );
  CIVX3 U923 ( .A(n915), .Z(n914) );
  CND2X4 U924 ( .A(n1972), .B(n2111), .Z(n915) );
  CNIVX1 U925 ( .A(n2303), .Z(n2338) );
  COND1XL U926 ( .A(n2398), .B(n2316), .C(n2380), .Z(\req_vec_rr_d[13][1] ) );
  CND3X1 U927 ( .A(n2383), .B(n2384), .C(n928), .Z(n2392) );
  CND3X2 U928 ( .A(n2164), .B(n2163), .C(n2162), .Z(n2165) );
  CND3X1 U929 ( .A(n2159), .B(n2158), .C(n2157), .Z(n2171) );
  CNIVX2 U930 ( .A(n2260), .Z(n2224) );
  CENXL U931 ( .A(n2313), .B(n2385), .Z(n2347) );
  CND2X1 U932 ( .A(n2154), .B(n2153), .Z(n2155) );
  COND1X2 U933 ( .A(n2239), .B(n2238), .C(n2237), .Z(n2259) );
  CIVX1 U934 ( .A(\req_vec_rr[3][2] ), .Z(n2232) );
  COND1X1 U935 ( .A(n2339), .B(n2338), .C(n2355), .Z(\req_vec_rr_d[1][2] ) );
  COND1X1 U936 ( .A(n2321), .B(n2338), .C(n2320), .Z(\req_vec_rr_d[15][0] ) );
  CIVX4 U937 ( .A(n2386), .Z(n2261) );
  CIVX3 U938 ( .A(n2224), .Z(n917) );
  COND1X1 U939 ( .A(n2319), .B(n2384), .C(n2383), .Z(\req_vec_rr_d[5][3] ) );
  CND2X2 U940 ( .A(n2384), .B(n2388), .Z(n2318) );
  CND2X4 U941 ( .A(n2384), .B(n2345), .Z(n2380) );
  CIVX8 U942 ( .A(n2385), .Z(n2361) );
  CANR1X2 U943 ( .A(\req_vec_rr[4][2] ), .B(n2286), .C(n2229), .Z(n2230) );
  CNR2IX2 U944 ( .B(n2328), .A(n1167), .Z(n1168) );
  CND2X4 U945 ( .A(n2037), .B(n2036), .Z(gnt_nxt[6]) );
  COR2XL U946 ( .A(n2224), .B(n2326), .Z(n928) );
  CNIVX3 U947 ( .A(n2326), .Z(n2320) );
  COR2XL U948 ( .A(n2326), .B(n2325), .Z(n978) );
  CNR3X2 U949 ( .A(n2279), .B(\req_vec_rr[15][0] ), .C(n2038), .Z(n1904) );
  CIVX4 U950 ( .A(n2260), .Z(n2345) );
  CND2X4 U951 ( .A(n2396), .B(n2365), .Z(n2367) );
  CNIVX1 U952 ( .A(\req_vec_rr[5][0] ), .Z(n918) );
  CNIVX1 U953 ( .A(\req_vec_rr[9][0] ), .Z(n919) );
  CNIVX1 U954 ( .A(\req_vec_rr[3][0] ), .Z(n920) );
  CNIVX1 U955 ( .A(\req_vec_rr[13][0] ), .Z(n921) );
  CNIVX1 U956 ( .A(\req_vec_rr[7][0] ), .Z(n922) );
  CNIVX1 U957 ( .A(\req_vec_rr[8][3] ), .Z(n923) );
  CNIVX1 U958 ( .A(\req_vec_rr[1][0] ), .Z(n924) );
  CNIVX1 U959 ( .A(n2404), .Z(n925) );
  CNIVX1 U960 ( .A(\req_vec_rr[6][1] ), .Z(n926) );
  COND1X1 U961 ( .A(n2295), .B(n2294), .C(n2293), .Z(n2296) );
  CND2X2 U962 ( .A(n2198), .B(n2197), .Z(n2201) );
  CND2X2 U963 ( .A(n2286), .B(\req_vec_rr[4][3] ), .Z(n2287) );
  CMXI2XL U964 ( .A0(n1398), .A1(n2394), .S(n2398), .Z(\req_vec_rr_d[5][2] )
         );
  CMXI2XL U965 ( .A0(n2379), .A1(n2378), .S(n2398), .Z(\req_vec_rr_d[9][3] )
         );
  CNIVX1 U966 ( .A(n1393), .Z(n927) );
  CNIVX12 U967 ( .A(req[3]), .Z(n1444) );
  CND2X2 U968 ( .A(n2358), .B(n2349), .Z(n2327) );
  CANR1X1 U969 ( .A(\req_vec_rr[1][0] ), .B(n2225), .C(n2146), .Z(n2149) );
  CIVDX2 U970 ( .A(n2191), .Z0(n1972), .Z1(n2146) );
  CNR2X2 U971 ( .A(n2396), .B(n934), .Z(n2310) );
  COR2X1 U972 ( .A(n1996), .B(n929), .Z(n930) );
  CIVX2 U973 ( .A(n1501), .Z(n929) );
  CND2X2 U974 ( .A(n2240), .B(n931), .Z(n1999) );
  CIVX20 U975 ( .A(n930), .Z(n931) );
  CND2X2 U976 ( .A(n1569), .B(n1570), .Z(n2215) );
  CND2X4 U977 ( .A(n2304), .B(n2389), .Z(n2306) );
  CND2X2 U978 ( .A(n1314), .B(n1287), .Z(n1265) );
  CANR1X2 U979 ( .A(n1731), .B(n1314), .C(n2328), .Z(n1128) );
  CNIVX1 U980 ( .A(n2375), .Z(n2394) );
  CNR2X2 U981 ( .A(n2297), .B(n2329), .Z(n1922) );
  CANR2X2 U982 ( .A(n1416), .B(n1717), .C(n1758), .D(n1421), .Z(n1208) );
  CANR1X2 U983 ( .A(n1976), .B(n1754), .C(n1691), .Z(n1693) );
  CNR2X4 U984 ( .A(n2154), .B(n2354), .Z(n1754) );
  CNR2IX4 U985 ( .B(n1502), .A(n2175), .Z(n2082) );
  CIVX4 U986 ( .A(n932), .Z(n934) );
  CNR2X4 U987 ( .A(n1578), .B(n1577), .Z(n1588) );
  CNR3X2 U988 ( .A(n2279), .B(\req_vec_rr[15][0] ), .C(n2079), .Z(n1970) );
  CNR3X2 U989 ( .A(n2279), .B(\req_vec_rr[15][0] ), .C(n1995), .Z(n1948) );
  CND2X2 U990 ( .A(n2147), .B(n1610), .Z(n1611) );
  CNR3X2 U991 ( .A(n2166), .B(\req_vec_rr[13][0] ), .C(\req_vec_rr[13][3] ), 
        .Z(n1502) );
  CNR2X2 U992 ( .A(n1012), .B(n1011), .Z(n1196) );
  CND3X2 U993 ( .A(n1004), .B(n1003), .C(n1002), .Z(n1005) );
  CANR1X2 U994 ( .A(n1153), .B(n1393), .C(\req_vec_rr[10][2] ), .Z(n1151) );
  CND3X1 U995 ( .A(n1058), .B(n1057), .C(n1072), .Z(n1059) );
  COND1X1 U996 ( .A(n1021), .B(n1419), .C(n1020), .Z(n1028) );
  CND2X1 U997 ( .A(n2225), .B(\req_vec_rr[1][2] ), .Z(n2226) );
  CNR2X2 U998 ( .A(n2060), .B(n2072), .Z(n2068) );
  CNIVX12 U999 ( .A(req[13]), .Z(n1428) );
  CND2X2 U1000 ( .A(n1428), .B(n1703), .Z(n1129) );
  CND4X2 U1001 ( .A(n2287), .B(n2289), .C(n2288), .D(n2290), .Z(n2295) );
  CND3X2 U1002 ( .A(n2204), .B(n1783), .C(n1954), .Z(n1180) );
  COND1X2 U1003 ( .A(n1975), .B(n1441), .C(n1303), .Z(n1305) );
  CNR2IX4 U1004 ( .B(n935), .A(n2261), .Z(n2375) );
  CIVX4 U1005 ( .A(n935), .Z(n2358) );
  CND4X2 U1006 ( .A(n1968), .B(n1967), .C(n1966), .D(n1965), .Z(n1969) );
  CNR2X4 U1007 ( .A(n2273), .B(\req_vec_rr[12][0] ), .Z(n1964) );
  COND1X2 U1008 ( .A(n2085), .B(n2084), .C(n2083), .Z(n2092) );
  CND3X4 U1009 ( .A(n1498), .B(n1497), .C(n1526), .Z(n2175) );
  CIVX3 U1010 ( .A(gnt_nxt[8]), .Z(n1994) );
  CND3X2 U1011 ( .A(n2270), .B(n1891), .C(n2322), .Z(n1894) );
  CND2X2 U1012 ( .A(n1113), .B(n1421), .Z(n1117) );
  CNIVX12 U1013 ( .A(req[11]), .Z(n1421) );
  COND1X2 U1014 ( .A(n1310), .B(n1421), .C(\req_vec_rr[1][3] ), .Z(n1311) );
  CANR1X2 U1015 ( .A(n1421), .B(n1443), .C(\req_vec_rr[2][2] ), .Z(n1422) );
  CND2X2 U1016 ( .A(n1155), .B(n1421), .Z(n1149) );
  CND2X2 U1017 ( .A(n1022), .B(n1421), .Z(n1026) );
  CND3X2 U1018 ( .A(n2204), .B(n1783), .C(n1736), .Z(n1640) );
  CND3X2 U1019 ( .A(n2204), .B(n2042), .C(n1954), .Z(n1895) );
  CNR2X1 U1020 ( .A(n2274), .B(n1890), .Z(n1898) );
  COR2X1 U1021 ( .A(n925), .B(n2384), .Z(n2393) );
  CND2X2 U1022 ( .A(n2313), .B(n2260), .Z(n935) );
  CNR2X4 U1023 ( .A(n1194), .B(n1195), .Z(n1199) );
  CND3X2 U1024 ( .A(n1016), .B(n1015), .C(n1014), .Z(n1017) );
  CND3X2 U1025 ( .A(n1009), .B(n1008), .C(n1007), .Z(n1012) );
  CIVXL U1026 ( .A(\req_vec_rr[14][2] ), .Z(n936) );
  CND2X1 U1027 ( .A(n1568), .B(n937), .Z(n2253) );
  CNR2X1 U1028 ( .A(n2173), .B(n936), .Z(n937) );
  CND3X4 U1029 ( .A(n1498), .B(n1497), .C(n1526), .Z(n938) );
  CND2X1 U1030 ( .A(n1023), .B(n1433), .Z(n1008) );
  CNR2X2 U1031 ( .A(n2171), .B(n2170), .Z(n2180) );
  CNR2X1 U1032 ( .A(n1872), .B(n2048), .Z(n1879) );
  CANR1X1 U1033 ( .A(n1408), .B(n1387), .C(n1386), .Z(n1390) );
  CANR2X1 U1034 ( .A(n1435), .B(n1084), .C(n1432), .D(n1085), .Z(n1082) );
  CND2X1 U1035 ( .A(n1393), .B(n1019), .Z(n1020) );
  COND1X1 U1036 ( .A(n1344), .B(n1343), .C(n1342), .Z(n1351) );
  COND1X2 U1037 ( .A(n1021), .B(n1343), .C(n1010), .Z(n1011) );
  CIVX2 U1038 ( .A(n2292), .Z(n2184) );
  CND2X1 U1039 ( .A(n1597), .B(n1596), .Z(n1599) );
  CNR3X1 U1040 ( .A(n2166), .B(\req_vec_rr[13][3] ), .C(n1889), .Z(n1573) );
  CNR2X2 U1041 ( .A(n2153), .B(\req_vec_rr[3][3] ), .Z(n1831) );
  CND2IX1 U1042 ( .B(n1189), .A(\req_vec_rr[15][3] ), .Z(n1098) );
  CIVX2 U1043 ( .A(n2151), .Z(n1847) );
  CNR2X1 U1044 ( .A(n1844), .B(n2023), .Z(n1837) );
  CND2X1 U1045 ( .A(n2236), .B(n2323), .Z(n2181) );
  CND2IX1 U1046 ( .B(n1870), .A(n2047), .Z(n1881) );
  COND1X1 U1047 ( .A(n1796), .B(n2110), .C(n1557), .Z(n1561) );
  CND3X1 U1048 ( .A(n2068), .B(n2067), .C(n2066), .Z(n2076) );
  CNR2X2 U1049 ( .A(n2046), .B(n2045), .Z(n2054) );
  CND3X1 U1050 ( .A(n1723), .B(n1722), .C(n1721), .Z(n1726) );
  CND2X1 U1051 ( .A(n1951), .B(n2005), .Z(n1946) );
  CND2IX1 U1052 ( .B(n1870), .A(n2005), .Z(n1822) );
  CND3X1 U1053 ( .A(n2031), .B(n2030), .C(n2029), .Z(n2034) );
  CND2X1 U1054 ( .A(n1762), .B(n2018), .Z(n1763) );
  CND3X1 U1055 ( .A(n1694), .B(n1693), .C(n1692), .Z(n1698) );
  CND2X1 U1056 ( .A(n1755), .B(n1971), .Z(n1694) );
  COND1XL U1057 ( .A(n2396), .B(n2322), .C(n2369), .Z(\req_vec_rr_d[10][0] )
         );
  CND2X1 U1058 ( .A(n2312), .B(n2318), .Z(\req_vec_rr_d[11][2] ) );
  CND2X2 U1059 ( .A(n2266), .B(n2265), .Z(n2324) );
  CANR3X1 U1060 ( .A(n1440), .B(n1087), .C(\req_vec_rr[13][2] ), .D(
        \req_vec_rr[13][3] ), .Z(n939) );
  CND2X1 U1061 ( .A(n1083), .B(n1400), .Z(n940) );
  CND3X2 U1062 ( .A(n940), .B(n1076), .C(n939), .Z(n1094) );
  CND2XL U1063 ( .A(n1371), .B(n1427), .Z(n941) );
  CANR1X1 U1064 ( .A(n1372), .B(n1363), .C(n1362), .Z(n942) );
  CND3X2 U1065 ( .A(n941), .B(n1364), .C(n942), .Z(n1382) );
  CNR2XL U1066 ( .A(n2026), .B(n1827), .Z(n943) );
  CND2X2 U1067 ( .A(n943), .B(n2147), .Z(n1828) );
  CND2IX1 U1068 ( .B(n2002), .A(n1874), .Z(n1816) );
  CND2XL U1069 ( .A(n2057), .B(n2113), .Z(n944) );
  CIVXL U1070 ( .A(n2058), .Z(n945) );
  COND2X1 U1071 ( .A(n2282), .B(n944), .C(n2116), .D(n945), .Z(n2060) );
  CND2IX2 U1072 ( .B(n2152), .A(n2319), .Z(n1853) );
  CND2XL U1073 ( .A(n2293), .B(n1971), .Z(n946) );
  COND1X1 U1074 ( .A(n1979), .B(n1978), .C(n2293), .Z(n947) );
  COND3X1 U1075 ( .A(n1981), .B(n946), .C(n1980), .D(n947), .Z(n1989) );
  CNR2XL U1076 ( .A(n1848), .B(n1798), .Z(n948) );
  CNR2X2 U1077 ( .A(n1807), .B(n948), .Z(n1800) );
  CND2IX1 U1078 ( .B(n1784), .A(n1874), .Z(n1785) );
  CND2IX1 U1079 ( .B(n2124), .A(n1757), .Z(n1690) );
  CNR2XL U1080 ( .A(\req_vec_rr[5][0] ), .B(\req_vec_rr[5][3] ), .Z(n949) );
  CND2X2 U1081 ( .A(n949), .B(n2283), .Z(n2110) );
  CND3XL U1082 ( .A(n1986), .B(n2114), .C(n2293), .Z(n950) );
  CND2XL U1083 ( .A(n1985), .B(n1984), .Z(n951) );
  CND3X1 U1084 ( .A(n951), .B(n1987), .C(n950), .Z(n1988) );
  CND2XL U1085 ( .A(n2352), .B(\req_vec_rr[6][2] ), .Z(n952) );
  CANR1X1 U1086 ( .A(n1372), .B(n1373), .C(n952), .Z(n1378) );
  CNR2X1 U1087 ( .A(n1031), .B(n1030), .Z(n953) );
  CND3XL U1088 ( .A(\req_vec_rr[15][3] ), .B(n1032), .C(n2317), .Z(n954) );
  COND2XL U1089 ( .A(n1419), .B(n1035), .C(n1034), .D(n1033), .Z(n955) );
  CND3XL U1090 ( .A(n1038), .B(n1036), .C(n1037), .Z(n956) );
  COND11X1 U1091 ( .A(n953), .B(n954), .C(n955), .D(n956), .Z(n1054) );
  CANR11X1 U1092 ( .A(\req_vec_rr[1][1] ), .B(\req_vec_rr[1][0] ), .C(n1314), 
        .D(n2339), .Z(n957) );
  CND2X1 U1093 ( .A(n1388), .B(n1315), .Z(n958) );
  CND4X2 U1094 ( .A(n1317), .B(n1316), .C(n957), .D(n958), .Z(n1318) );
  CND2IX1 U1095 ( .B(n2090), .A(n1874), .Z(n1583) );
  CND2X1 U1096 ( .A(n1850), .B(n1799), .Z(n959) );
  CND2X1 U1097 ( .A(n959), .B(n1800), .Z(n960) );
  CANR1X2 U1098 ( .A(n1831), .B(n1801), .C(n960), .Z(n1806) );
  CND2X1 U1099 ( .A(n1825), .B(n2018), .Z(n961) );
  COND1X1 U1100 ( .A(n2017), .B(n1853), .C(n961), .Z(n1841) );
  CND2IXL U1101 ( .B(n1621), .A(n2236), .Z(n1622) );
  CND2IXL U1102 ( .B(n2032), .A(n2146), .Z(n2033) );
  CNR2IX1 U1103 ( .B(n1428), .A(n1245), .Z(n1249) );
  CNR2XL U1104 ( .A(\req_vec_rr[1][0] ), .B(n2374), .Z(n962) );
  CND2X1 U1105 ( .A(n1384), .B(n962), .Z(n1316) );
  CANR1X1 U1106 ( .A(n1433), .B(n1087), .C(n1081), .Z(n963) );
  CND2XL U1107 ( .A(n1083), .B(n1434), .Z(n964) );
  CND3X2 U1108 ( .A(n964), .B(n1082), .C(n963), .Z(n1092) );
  CNR2XL U1109 ( .A(\req_vec_rr[8][3] ), .B(n2314), .Z(n965) );
  CND2X1 U1110 ( .A(n2247), .B(n965), .Z(n2089) );
  CNR3X2 U1111 ( .A(n1614), .B(n1615), .C(n2334), .Z(n966) );
  CND2X2 U1112 ( .A(n1616), .B(n966), .Z(n2151) );
  CND2IXL U1113 ( .B(n2026), .A(n1757), .Z(n1761) );
  CND2X1 U1114 ( .A(n2326), .B(n2325), .Z(n967) );
  CND2X2 U1115 ( .A(n967), .B(n2386), .Z(n2353) );
  CND2IXL U1116 ( .B(n1807), .A(n2236), .Z(n1808) );
  CNR2X1 U1117 ( .A(n2121), .B(n2129), .Z(n968) );
  CND2X1 U1118 ( .A(n2112), .B(n2111), .Z(n969) );
  CND3X1 U1119 ( .A(n969), .B(n968), .C(n2128), .Z(n2131) );
  CIVXL U1120 ( .A(\req_vec_rr[3][2] ), .Z(n970) );
  COND1XL U1121 ( .A(n2398), .B(n970), .C(n2318), .Z(\req_vec_rr_d[3][2] ) );
  CIVXL U1122 ( .A(\req_vec_rr[4][0] ), .Z(n971) );
  COND1X1 U1123 ( .A(n971), .B(n2356), .C(n2369), .Z(\req_vec_rr_d[4][0] ) );
  CND2IX1 U1124 ( .B(\req_vec_rr[3][2] ), .A(\req_vec_rr[3][3] ), .Z(n1321) );
  CNR2IX1 U1125 ( .B(n1433), .A(n1245), .Z(n1227) );
  CND2IX1 U1126 ( .B(n2166), .A(\req_vec_rr[13][3] ), .Z(n1183) );
  CNR2IX1 U1127 ( .B(n2069), .A(\req_vec_rr[6][3] ), .Z(n1846) );
  CND2IX1 U1128 ( .B(n2353), .A(n2327), .Z(n2370) );
  CND2IX1 U1129 ( .B(n1837), .A(n1838), .Z(n1839) );
  CND2IX1 U1130 ( .B(n2129), .A(n2199), .Z(n2130) );
  CND2X1 U1131 ( .A(n2365), .B(\req_vec_rr[2][1] ), .Z(n972) );
  CND2X1 U1132 ( .A(n2367), .B(n972), .Z(\req_vec_rr_d[2][1] ) );
  COAN1X1 U1133 ( .A(n924), .B(n2384), .C(n2369), .Z(n2405) );
  CIVX4 U1134 ( .A(\req_vec_rr[5][3] ), .Z(n2319) );
  CAN3X2 U1135 ( .A(n1331), .B(n1330), .C(n1329), .Z(n973) );
  COAN1X2 U1136 ( .A(n1424), .B(n1419), .C(n1418), .Z(n974) );
  CAN2X1 U1137 ( .A(n1441), .B(n1376), .Z(n975) );
  CAN2X1 U1138 ( .A(n1753), .B(n2015), .Z(n976) );
  CAN4X1 U1139 ( .A(n2275), .B(n2274), .C(n2273), .D(n2272), .Z(n977) );
  CIVDX2 U1140 ( .A(n1695), .Z0(n1982), .Z1(n2199) );
  CIVDX3 U1141 ( .A(n1695), .Z0(n2293), .Z1(n2236) );
  CIVX4 U1142 ( .A(\req_vec_rr[8][2] ), .Z(n2328) );
  CAN2X1 U1143 ( .A(n1736), .B(n2042), .Z(n979) );
  COR2XL U1144 ( .A(n1774), .B(\req_vec_rr[15][0] ), .Z(n980) );
  CMXI2XL U1145 ( .A0(n2371), .A1(n2385), .S(n2398), .Z(\req_vec_rr_d[7][3] )
         );
  CND2X2 U1146 ( .A(n1612), .B(n1611), .Z(n1613) );
  CND2X4 U1147 ( .A(n2211), .B(n2280), .Z(n2222) );
  CND3X2 U1148 ( .A(n2204), .B(n2000), .C(n1954), .Z(n1938) );
  CND2X2 U1149 ( .A(n2281), .B(n2280), .Z(n2298) );
  CIVX3 U1150 ( .A(n1175), .Z(n1177) );
  CND2XL U1151 ( .A(n1936), .B(n1731), .Z(n1739) );
  CND2X1 U1152 ( .A(n1936), .B(n1703), .Z(n1638) );
  CNR2X2 U1153 ( .A(n1435), .B(n1798), .Z(n1307) );
  CIVX2 U1154 ( .A(n1522), .Z(n1192) );
  CNIVX8 U1157 ( .A(req[2]), .Z(n1441) );
  CNR2IX1 U1158 ( .B(\req_vec_rr[12][1] ), .A(\req_vec_rr[12][0] ), .Z(n995)
         );
  CNR2X1 U1159 ( .A(\req_vec_rr[12][1] ), .B(\req_vec_rr[12][0] ), .Z(n994) );
  CIVX3 U1160 ( .A(req[0]), .Z(n981) );
  CIVX8 U1161 ( .A(n981), .Z(n1445) );
  CANR2X1 U1162 ( .A(n1441), .B(n995), .C(n994), .D(n1445), .Z(n984) );
  CNIVX8 U1163 ( .A(req[1]), .Z(n1440) );
  CNR2IX2 U1164 ( .B(\req_vec_rr[12][0] ), .A(\req_vec_rr[12][1] ), .Z(n996)
         );
  CANR3X1 U1165 ( .A(n1440), .B(n996), .C(\req_vec_rr[12][3] ), .D(
        \req_vec_rr[12][2] ), .Z(n983) );
  CAN2X1 U1166 ( .A(\req_vec_rr[12][1] ), .B(\req_vec_rr[12][0] ), .Z(n997) );
  CND2X1 U1167 ( .A(n1444), .B(n997), .Z(n982) );
  CND3X2 U1168 ( .A(n984), .B(n983), .C(n982), .Z(n1494) );
  CNIVX4 U1169 ( .A(req[14]), .Z(n1384) );
  CIVX3 U1170 ( .A(req[12]), .Z(n985) );
  CIVX8 U1171 ( .A(n985), .Z(n1388) );
  CANR2X1 U1172 ( .A(n1384), .B(n995), .C(n994), .D(n1388), .Z(n989) );
  CND2X1 U1173 ( .A(\req_vec_rr[12][2] ), .B(\req_vec_rr[12][3] ), .Z(n986) );
  CANR1X1 U1174 ( .A(n996), .B(n1428), .C(n986), .Z(n988) );
  CNIVX4 U1175 ( .A(req[15]), .Z(n1426) );
  CND2X1 U1176 ( .A(n1426), .B(n997), .Z(n987) );
  CND3X2 U1177 ( .A(n989), .B(n988), .C(n987), .Z(n1493) );
  CNIVX8 U1178 ( .A(req[10]), .Z(n1392) );
  CIVX3 U1179 ( .A(req[8]), .Z(n990) );
  CIVX8 U1180 ( .A(n990), .Z(n1393) );
  CANR2X1 U1181 ( .A(n1392), .B(n995), .C(n994), .D(n1393), .Z(n993) );
  CNIVX8 U1182 ( .A(req[9]), .Z(n1416) );
  CANR3X2 U1183 ( .A(n996), .B(n1416), .C(n2413), .D(\req_vec_rr[12][2] ), .Z(
        n992) );
  CND2X1 U1184 ( .A(n1421), .B(n997), .Z(n991) );
  CND3X2 U1185 ( .A(n993), .B(n992), .C(n991), .Z(n1492) );
  CNIVX8 U1186 ( .A(req[6]), .Z(n1432) );
  CNIVX4 U1187 ( .A(req[4]), .Z(n1341) );
  CANR2X1 U1188 ( .A(n1432), .B(n995), .C(n994), .D(n1341), .Z(n1000) );
  CNIVX16 U1189 ( .A(req[5]), .Z(n1433) );
  CIVX2 U1190 ( .A(\req_vec_rr[12][2] ), .Z(n2243) );
  CANR3X2 U1191 ( .A(n996), .B(n1433), .C(n2243), .D(\req_vec_rr[12][3] ), .Z(
        n999) );
  CNIVX16 U1192 ( .A(req[7]), .Z(n1434) );
  CND2X1 U1193 ( .A(n1434), .B(n997), .Z(n998) );
  CND3X2 U1194 ( .A(n1000), .B(n999), .C(n998), .Z(n1491) );
  CND4X2 U1195 ( .A(n1494), .B(n1493), .C(n1492), .D(n1491), .Z(n1524) );
  CIVX4 U1196 ( .A(\req_vec_rr[11][0] ), .Z(n1635) );
  CND2X1 U1197 ( .A(n1635), .B(\req_vec_rr[11][1] ), .Z(n1021) );
  CNR2X2 U1198 ( .A(\req_vec_rr[11][0] ), .B(\req_vec_rr[11][1] ), .Z(n1019)
         );
  CND2X1 U1199 ( .A(n1019), .B(n1445), .Z(n1001) );
  COND1X2 U1200 ( .A(n1021), .B(n1334), .C(n1001), .Z(n1006) );
  CIVX2 U1201 ( .A(\req_vec_rr[11][1] ), .Z(n2342) );
  CNR2X2 U1202 ( .A(n2342), .B(n1635), .Z(n1022) );
  CND2X1 U1203 ( .A(n1022), .B(n1444), .Z(n1004) );
  CNR2X2 U1204 ( .A(n1635), .B(\req_vec_rr[11][1] ), .Z(n1023) );
  CND2X1 U1205 ( .A(n1023), .B(n1440), .Z(n1003) );
  CNR2X1 U1206 ( .A(\req_vec_rr[11][3] ), .B(\req_vec_rr[11][2] ), .Z(n1002)
         );
  CNR2X2 U1207 ( .A(n1006), .B(n1005), .Z(n1197) );
  CND2X1 U1208 ( .A(n1022), .B(n1434), .Z(n1009) );
  CIVDX1 U1209 ( .A(\req_vec_rr[11][2] ), .Z0(n1580) );
  CNR2X1 U1210 ( .A(\req_vec_rr[11][3] ), .B(n1580), .Z(n1007) );
  CIVX4 U1211 ( .A(n1432), .Z(n1343) );
  CND2X2 U1212 ( .A(n1341), .B(n1019), .Z(n1010) );
  CNR2X2 U1213 ( .A(n1197), .B(n1196), .Z(n1029) );
  CNIVX4 U1214 ( .A(req[14]), .Z(n1425) );
  CIVX2 U1215 ( .A(n1425), .Z(n1246) );
  CND2X1 U1216 ( .A(n1019), .B(n1388), .Z(n1013) );
  COND1X1 U1217 ( .A(n1021), .B(n1246), .C(n1013), .Z(n1018) );
  CND2X1 U1218 ( .A(n1023), .B(n1428), .Z(n1016) );
  CND2X1 U1219 ( .A(n1426), .B(n1022), .Z(n1015) );
  CIVX2 U1220 ( .A(\req_vec_rr[11][3] ), .Z(n1634) );
  CNR2X1 U1221 ( .A(n1634), .B(n1580), .Z(n1014) );
  CNR2X2 U1222 ( .A(n1018), .B(n1017), .Z(n1195) );
  CIVX8 U1223 ( .A(n1392), .Z(n1419) );
  CND2X1 U1224 ( .A(n1023), .B(n1416), .Z(n1025) );
  CNR2X1 U1225 ( .A(n1634), .B(\req_vec_rr[11][2] ), .Z(n1024) );
  CND3X2 U1226 ( .A(n1026), .B(n1025), .C(n1024), .Z(n1027) );
  CNR2X2 U1227 ( .A(n1028), .B(n1027), .Z(n1194) );
  CND2X4 U1228 ( .A(n1029), .B(n1199), .Z(n1629) );
  CND2X2 U1229 ( .A(n1629), .B(n1524), .Z(n1189) );
  CNIVX4 U1230 ( .A(n1416), .Z(n1240) );
  CIVXL U1231 ( .A(n1240), .Z(n1031) );
  CIVX2 U1232 ( .A(\req_vec_rr[15][0] ), .Z(n2321) );
  CNR2X1 U1233 ( .A(n2321), .B(\req_vec_rr[15][1] ), .Z(n1047) );
  CIVX1 U1234 ( .A(n1047), .Z(n1030) );
  CNR2X1 U1235 ( .A(\req_vec_rr[15][1] ), .B(\req_vec_rr[15][0] ), .Z(n1043)
         );
  CNIVX4 U1236 ( .A(n1393), .Z(n1420) );
  CND2X1 U1237 ( .A(n1043), .B(n1420), .Z(n1032) );
  CIVX2 U1238 ( .A(\req_vec_rr[15][2] ), .Z(n2317) );
  CIVX2 U1239 ( .A(\req_vec_rr[15][1] ), .Z(n2337) );
  CNR2X1 U1240 ( .A(n2337), .B(\req_vec_rr[15][0] ), .Z(n1044) );
  CIVX1 U1241 ( .A(n1044), .Z(n1035) );
  CIVX2 U1242 ( .A(n1421), .Z(n1034) );
  CNR2X1 U1243 ( .A(n2337), .B(n2321), .Z(n1046) );
  CIVX1 U1244 ( .A(n1046), .Z(n1033) );
  CANR3XL U1245 ( .A(n1046), .B(n1444), .C(\req_vec_rr[15][3] ), .D(
        \req_vec_rr[15][2] ), .Z(n1038) );
  CIVDX2 U1246 ( .A(n1441), .Z0(n1334), .Z1(n1222) );
  CIVX2 U1247 ( .A(n1445), .Z(n1218) );
  CIVX2 U1248 ( .A(n1218), .Z(n1366) );
  CANR2X1 U1249 ( .A(n1044), .B(n1222), .C(n1366), .D(n1043), .Z(n1037) );
  CNIVX4 U1250 ( .A(n1440), .Z(n1365) );
  CND2X1 U1251 ( .A(n1047), .B(n1365), .Z(n1036) );
  CNIVX2 U1252 ( .A(n1432), .Z(n1375) );
  CNIVX4 U1253 ( .A(req[4]), .Z(n1435) );
  CNIVX4 U1254 ( .A(n1435), .Z(n1370) );
  CANR2X1 U1255 ( .A(n1044), .B(n1375), .C(n1370), .D(n1043), .Z(n1042) );
  CNIVX4 U1256 ( .A(n1434), .Z(n1373) );
  CND2XL U1257 ( .A(n1046), .B(n1373), .Z(n1041) );
  CND2X1 U1258 ( .A(n1047), .B(n1433), .Z(n1040) );
  CNR2X1 U1259 ( .A(n2317), .B(\req_vec_rr[15][3] ), .Z(n1039) );
  CND4X1 U1260 ( .A(n1042), .B(n1041), .C(n1040), .D(n1039), .Z(n1052) );
  CNIVX4 U1261 ( .A(n1384), .Z(n1361) );
  CNIVX4 U1262 ( .A(n1388), .Z(n1427) );
  CANR2XL U1263 ( .A(n1044), .B(n1361), .C(n1427), .D(n1043), .Z(n1050) );
  CNIVX4 U1264 ( .A(n1426), .Z(n1363) );
  CND2X1 U1265 ( .A(\req_vec_rr[15][3] ), .B(\req_vec_rr[15][2] ), .Z(n1045)
         );
  CANR1XL U1266 ( .A(n1363), .B(n1046), .C(n1045), .Z(n1049) );
  CNIVX4 U1267 ( .A(n1428), .Z(n1360) );
  CND2XL U1268 ( .A(n1047), .B(n1360), .Z(n1048) );
  CND3X1 U1269 ( .A(n1050), .B(n1049), .C(n1048), .Z(n1051) );
  CND2X1 U1270 ( .A(n1052), .B(n1051), .Z(n1053) );
  CNR2X2 U1271 ( .A(n1054), .B(n1053), .Z(n1097) );
  CIVX2 U1272 ( .A(\req_vec_rr[14][1] ), .Z(n1743) );
  CIVX4 U1273 ( .A(\req_vec_rr[14][0] ), .Z(n2183) );
  CNR2X1 U1274 ( .A(n1743), .B(n2183), .Z(n1067) );
  CNR2X2 U1275 ( .A(\req_vec_rr[14][1] ), .B(\req_vec_rr[14][0] ), .Z(n1066)
         );
  CANR2X1 U1276 ( .A(n1067), .B(n1363), .C(n1388), .D(n1066), .Z(n1056) );
  CNR2X2 U1277 ( .A(n1743), .B(\req_vec_rr[14][0] ), .Z(n1065) );
  CNR2X2 U1278 ( .A(\req_vec_rr[14][1] ), .B(n2183), .Z(n1064) );
  CANR2X2 U1279 ( .A(n1065), .B(n1361), .C(n1428), .D(n1064), .Z(n1055) );
  CND3X2 U1280 ( .A(n1056), .B(n1055), .C(\req_vec_rr[14][2] ), .Z(n1060) );
  CANR2X1 U1281 ( .A(n1067), .B(n1421), .C(n1066), .D(n1393), .Z(n1058) );
  CANR2X1 U1282 ( .A(n1065), .B(n1392), .C(n1416), .D(n1064), .Z(n1057) );
  CND2X2 U1283 ( .A(n1060), .B(n1059), .Z(n1061) );
  CND2IX2 U1284 ( .B(n2404), .A(n1061), .Z(n1075) );
  CIVX2 U1285 ( .A(\req_vec_rr[14][2] ), .Z(n1072) );
  CANR2X1 U1286 ( .A(n1067), .B(n1434), .C(n1435), .D(n1066), .Z(n1063) );
  CANR2X1 U1287 ( .A(n1064), .B(n1433), .C(n1065), .D(n1432), .Z(n1062) );
  CND2X1 U1288 ( .A(n1063), .B(n1062), .Z(n1071) );
  CANR2X1 U1289 ( .A(n1065), .B(n1441), .C(n1440), .D(n1064), .Z(n1069) );
  CANR2X1 U1290 ( .A(n1067), .B(n1444), .C(n1445), .D(n1066), .Z(n1068) );
  CND3X2 U1291 ( .A(n1069), .B(n1068), .C(n1072), .Z(n1070) );
  COND1X2 U1292 ( .A(n1072), .B(n1071), .C(n1070), .Z(n1073) );
  CND2IX2 U1293 ( .B(n2403), .A(n1073), .Z(n1074) );
  CND2X4 U1294 ( .A(n1075), .B(n1074), .Z(n1522) );
  CIVX4 U1295 ( .A(\req_vec_rr[13][0] ), .Z(n1889) );
  CNR2X2 U1296 ( .A(n1889), .B(\req_vec_rr[13][1] ), .Z(n1087) );
  CIVX2 U1297 ( .A(\req_vec_rr[13][1] ), .Z(n2316) );
  CNR2X2 U1298 ( .A(n1889), .B(n2316), .Z(n1083) );
  CNIVX4 U1299 ( .A(n1444), .Z(n1400) );
  CNR2X1 U1300 ( .A(\req_vec_rr[13][0] ), .B(\req_vec_rr[13][1] ), .Z(n1084)
         );
  CNR2IX1 U1301 ( .B(\req_vec_rr[13][1] ), .A(\req_vec_rr[13][0] ), .Z(n1085)
         );
  CANR2X1 U1302 ( .A(n1445), .B(n1084), .C(n1441), .D(n1085), .Z(n1076) );
  CANR2X1 U1303 ( .A(n1085), .B(n1392), .C(n1084), .D(n1393), .Z(n1080) );
  CND2IX1 U1304 ( .B(\req_vec_rr[13][2] ), .A(\req_vec_rr[13][3] ), .Z(n1077)
         );
  CANR1X1 U1305 ( .A(n1416), .B(n1087), .C(n1077), .Z(n1079) );
  CND2X1 U1306 ( .A(n1083), .B(n1421), .Z(n1078) );
  CND3X1 U1307 ( .A(n1080), .B(n1079), .C(n1078), .Z(n1093) );
  CND2IX1 U1308 ( .B(\req_vec_rr[13][3] ), .A(\req_vec_rr[13][2] ), .Z(n1081)
         );
  CND2X1 U1309 ( .A(n1083), .B(n1363), .Z(n1090) );
  CANR2X1 U1310 ( .A(n1384), .B(n1085), .C(n1084), .D(n1388), .Z(n1089) );
  CND2X1 U1311 ( .A(\req_vec_rr[13][2] ), .B(\req_vec_rr[13][3] ), .Z(n1086)
         );
  CANR1X1 U1312 ( .A(n1428), .B(n1087), .C(n1086), .Z(n1088) );
  CND3X2 U1313 ( .A(n1090), .B(n1089), .C(n1088), .Z(n1091) );
  CND4X4 U1314 ( .A(n1094), .B(n1093), .C(n1092), .D(n1091), .Z(n2166) );
  CND2X2 U1315 ( .A(n1522), .B(n2166), .Z(n1095) );
  CIVX3 U1316 ( .A(n1095), .Z(n1096) );
  CND2X4 U1317 ( .A(n1097), .B(n1096), .Z(n2174) );
  CNR2X4 U1318 ( .A(n1098), .B(n2174), .Z(n1627) );
  CNR2IX2 U1319 ( .B(\req_vec_rr[9][1] ), .A(\req_vec_rr[9][0] ), .Z(n1112) );
  CNR2X1 U1320 ( .A(\req_vec_rr[9][0] ), .B(\req_vec_rr[9][1] ), .Z(n1111) );
  CANR2X2 U1321 ( .A(n1112), .B(n1441), .C(n1111), .D(n1445), .Z(n1101) );
  CIVX3 U1322 ( .A(\req_vec_rr[9][0] ), .Z(n1628) );
  CNIVX4 U1323 ( .A(\req_vec_rr[9][1] ), .Z(n2203) );
  CNR2X2 U1324 ( .A(n1628), .B(n2203), .Z(n1115) );
  CANR3X2 U1325 ( .A(n1115), .B(n1440), .C(\req_vec_rr[9][2] ), .D(
        \req_vec_rr[9][3] ), .Z(n1100) );
  CIVX2 U1326 ( .A(\req_vec_rr[9][1] ), .Z(n2381) );
  CNR2X2 U1327 ( .A(n1628), .B(n2381), .Z(n1113) );
  CND2X1 U1328 ( .A(n1113), .B(n1444), .Z(n1099) );
  CND3X2 U1329 ( .A(n1101), .B(n1100), .C(n1099), .Z(n1122) );
  CANR2X2 U1330 ( .A(n1111), .B(n1435), .C(n1112), .D(n1432), .Z(n1105) );
  CND2IX1 U1331 ( .B(\req_vec_rr[9][3] ), .A(\req_vec_rr[9][2] ), .Z(n1102) );
  CANR1X1 U1332 ( .A(n1433), .B(n1115), .C(n1102), .Z(n1104) );
  CND2X1 U1333 ( .A(n1113), .B(n1434), .Z(n1103) );
  CND3X2 U1334 ( .A(n1105), .B(n1104), .C(n1103), .Z(n1121) );
  CND2X1 U1335 ( .A(\req_vec_rr[9][3] ), .B(\req_vec_rr[9][2] ), .Z(n1106) );
  CANR1X1 U1336 ( .A(n1113), .B(n1426), .C(n1106), .Z(n1110) );
  CND2X1 U1337 ( .A(n1388), .B(n1111), .Z(n1109) );
  CND2X2 U1338 ( .A(n1428), .B(n1115), .Z(n1108) );
  CND2X1 U1339 ( .A(n1425), .B(n1112), .Z(n1107) );
  CND4X2 U1340 ( .A(n1110), .B(n1109), .C(n1108), .D(n1107), .Z(n1120) );
  CANR2X2 U1341 ( .A(n1112), .B(n1392), .C(n1111), .D(n1393), .Z(n1118) );
  CIVX2 U1342 ( .A(\req_vec_rr[9][2] ), .Z(n2357) );
  CND2X1 U1343 ( .A(\req_vec_rr[9][3] ), .B(n2357), .Z(n1114) );
  CANR1X2 U1344 ( .A(n1115), .B(n1416), .C(n1114), .Z(n1116) );
  CND3X2 U1345 ( .A(n1118), .B(n1117), .C(n1116), .Z(n1119) );
  CND4X4 U1346 ( .A(n1122), .B(n1121), .C(n1120), .D(n1119), .Z(n1173) );
  CNIVX4 U1347 ( .A(\req_vec_rr[8][0] ), .Z(n2314) );
  CNR2X4 U1348 ( .A(n2314), .B(\req_vec_rr[8][1] ), .Z(n1892) );
  CANR1X1 U1349 ( .A(n1892), .B(n1393), .C(\req_vec_rr[8][2] ), .Z(n1126) );
  CAN2X2 U1350 ( .A(\req_vec_rr[8][0] ), .B(\req_vec_rr[8][1] ), .Z(n1731) );
  CND2X1 U1351 ( .A(n1421), .B(n1731), .Z(n1125) );
  CNR2IX2 U1352 ( .B(\req_vec_rr[8][1] ), .A(\req_vec_rr[8][0] ), .Z(n1955) );
  CND2X1 U1353 ( .A(n1392), .B(n1955), .Z(n1124) );
  CNR2IX2 U1354 ( .B(\req_vec_rr[8][0] ), .A(\req_vec_rr[8][1] ), .Z(n1703) );
  CND2X1 U1355 ( .A(n1416), .B(n1703), .Z(n1123) );
  CND4X2 U1356 ( .A(n1126), .B(n1125), .C(n1124), .D(n1123), .Z(n1165) );
  CNIVX2 U1357 ( .A(req[15]), .Z(n1314) );
  CANR2X2 U1358 ( .A(n1955), .B(n1384), .C(n1892), .D(n1388), .Z(n1127) );
  CANR11X4 U1359 ( .A(n1129), .B(n1128), .C(n1127), .D(n2414), .Z(n1164) );
  CND2X4 U1360 ( .A(n1165), .B(n1164), .Z(n1676) );
  CNR2IX2 U1361 ( .B(\req_vec_rr[10][0] ), .A(\req_vec_rr[10][1] ), .Z(n1152)
         );
  CIVX2 U1362 ( .A(\req_vec_rr[10][1] ), .Z(n2216) );
  CIVX2 U1363 ( .A(\req_vec_rr[10][0] ), .Z(n2322) );
  CNR2X2 U1364 ( .A(n2216), .B(n2322), .Z(n1155) );
  CANR2X2 U1365 ( .A(n1152), .B(n1433), .C(n1155), .D(n1434), .Z(n1132) );
  CNR2X2 U1366 ( .A(\req_vec_rr[10][1] ), .B(\req_vec_rr[10][0] ), .Z(n1153)
         );
  CND2X1 U1367 ( .A(n1153), .B(n1435), .Z(n1131) );
  CNR2X2 U1368 ( .A(n2216), .B(\req_vec_rr[10][0] ), .Z(n1154) );
  CIVX2 U1369 ( .A(\req_vec_rr[10][2] ), .Z(n2262) );
  CANR1X1 U1370 ( .A(n1432), .B(n1154), .C(n2262), .Z(n1130) );
  CND3X2 U1371 ( .A(n1132), .B(n1131), .C(n1130), .Z(n1137) );
  CANR2X2 U1372 ( .A(n1154), .B(n1441), .C(n1445), .D(n1153), .Z(n1135) );
  CANR1X1 U1373 ( .A(n1444), .B(n1155), .C(\req_vec_rr[10][2] ), .Z(n1134) );
  CND2X1 U1374 ( .A(n1152), .B(n1440), .Z(n1133) );
  CND3X2 U1375 ( .A(n1135), .B(n1134), .C(n1133), .Z(n1136) );
  CND3X4 U1376 ( .A(n1137), .B(n1136), .C(n2416), .Z(n1489) );
  CND3X2 U1377 ( .A(n1173), .B(n1676), .C(n1489), .Z(n1184) );
  CND2X2 U1378 ( .A(n1432), .B(n1955), .Z(n1505) );
  CIVX3 U1379 ( .A(n1505), .Z(n1139) );
  CND2X2 U1380 ( .A(n1341), .B(n1892), .Z(n1507) );
  CIVX3 U1381 ( .A(n1507), .Z(n1138) );
  CNR2X4 U1382 ( .A(n1139), .B(n1138), .Z(n1142) );
  CND2X4 U1383 ( .A(n1433), .B(n1703), .Z(n1508) );
  CND2X4 U1384 ( .A(n1434), .B(n1731), .Z(n1504) );
  CND3X4 U1385 ( .A(n1508), .B(n1504), .C(\req_vec_rr[8][2] ), .Z(n1140) );
  CIVX4 U1386 ( .A(n1140), .Z(n1141) );
  CND2X4 U1387 ( .A(n1142), .B(n1141), .Z(n1171) );
  CND2X2 U1388 ( .A(n1440), .B(n1703), .Z(n1144) );
  CND2X2 U1389 ( .A(n1441), .B(n1955), .Z(n1143) );
  CND2X4 U1390 ( .A(n1144), .B(n1143), .Z(n1166) );
  CND2X2 U1391 ( .A(n1445), .B(n1892), .Z(n1146) );
  CND2X4 U1392 ( .A(n1444), .B(n1731), .Z(n1145) );
  CND2X4 U1393 ( .A(n1146), .B(n1145), .Z(n1167) );
  CNR2X2 U1394 ( .A(n1166), .B(n1167), .Z(n1513) );
  CND2X2 U1395 ( .A(n1513), .B(n2328), .Z(n1147) );
  CND3X2 U1396 ( .A(n1171), .B(n1147), .C(n2414), .Z(n1161) );
  CND2X1 U1397 ( .A(n1154), .B(n1392), .Z(n1150) );
  CND2X1 U1398 ( .A(n1152), .B(n1416), .Z(n1148) );
  CND4X1 U1399 ( .A(n1151), .B(n1150), .C(n1149), .D(n1148), .Z(n1160) );
  CANR2X2 U1400 ( .A(n1388), .B(n1153), .C(n1152), .D(n1428), .Z(n1158) );
  CANR1X1 U1401 ( .A(n1384), .B(n1154), .C(n2262), .Z(n1157) );
  CND2X1 U1402 ( .A(n1426), .B(n1155), .Z(n1156) );
  CND3X2 U1403 ( .A(n1158), .B(n1157), .C(n1156), .Z(n1159) );
  CND3X4 U1404 ( .A(n1160), .B(n1159), .C(\req_vec_rr[10][3] ), .Z(n1490) );
  CND2X4 U1405 ( .A(n1161), .B(n1490), .Z(n1529) );
  CNR2X4 U1406 ( .A(n1184), .B(n1529), .Z(n2144) );
  CIVX4 U1407 ( .A(n2144), .Z(n1643) );
  CIVX8 U1408 ( .A(n1643), .Z(n2276) );
  CND2X4 U1409 ( .A(n1627), .B(n2276), .Z(n2279) );
  CND2X1 U1410 ( .A(n2337), .B(\req_vec_rr[15][2] ), .Z(n1774) );
  CNR2X1 U1411 ( .A(n2279), .B(n980), .Z(n1456) );
  CAN3X2 U1412 ( .A(n1173), .B(n1676), .C(n1489), .Z(n1631) );
  CND2XL U1413 ( .A(n1635), .B(\req_vec_rr[11][3] ), .Z(n1162) );
  CNR3X1 U1414 ( .A(n1529), .B(n1629), .C(n1162), .Z(n1163) );
  CND2X1 U1415 ( .A(n1631), .B(n1163), .Z(n1952) );
  CNR2X1 U1416 ( .A(\req_vec_rr[11][1] ), .B(n1580), .Z(n1636) );
  CIVX2 U1417 ( .A(n1636), .Z(n1782) );
  CNR2X1 U1418 ( .A(n1952), .B(n1782), .Z(n1182) );
  CIVX2 U1419 ( .A(n1173), .Z(n1172) );
  CND2X4 U1420 ( .A(n1165), .B(n1164), .Z(n1516) );
  CIVX3 U1421 ( .A(n1166), .Z(n1169) );
  CND2X4 U1422 ( .A(n1169), .B(n1168), .Z(n1170) );
  CND3X4 U1423 ( .A(n1171), .B(n1170), .C(n2414), .Z(n1174) );
  CND3X4 U1424 ( .A(n1172), .B(n1516), .C(n1174), .Z(n2268) );
  CIVX8 U1425 ( .A(n2268), .Z(n2204) );
  CNR2IX1 U1426 ( .B(\req_vec_rr[9][2] ), .A(n2203), .Z(n1783) );
  CIVX2 U1427 ( .A(\req_vec_rr[9][3] ), .Z(n2379) );
  CNR2X1 U1428 ( .A(n2379), .B(\req_vec_rr[9][0] ), .Z(n1954) );
  CND2X4 U1429 ( .A(n1174), .B(n1173), .Z(n1500) );
  CIVX2 U1430 ( .A(n1500), .Z(n1175) );
  CND2IX1 U1431 ( .B(n1490), .A(n1516), .Z(n1176) );
  CNR2X4 U1432 ( .A(n1177), .B(n1176), .Z(n2270) );
  CNR2X1 U1433 ( .A(\req_vec_rr[10][1] ), .B(n2262), .Z(n1642) );
  CND3X1 U1434 ( .A(n2270), .B(n2322), .C(n1642), .Z(n1179) );
  CNR2X1 U1435 ( .A(n1516), .B(n2328), .Z(n1936) );
  CND2X1 U1436 ( .A(n1936), .B(n1892), .Z(n1178) );
  CND3X2 U1437 ( .A(n1179), .B(n1180), .C(n1178), .Z(n1181) );
  CNR2X2 U1438 ( .A(n1182), .B(n1181), .Z(n1204) );
  CNR2X2 U1439 ( .A(n1189), .B(n1183), .Z(n1188) );
  CNIVX1 U1440 ( .A(n1184), .Z(n1185) );
  CIVX2 U1441 ( .A(n1185), .Z(n1187) );
  CNIVX4 U1442 ( .A(n1529), .Z(n1632) );
  CIVX3 U1443 ( .A(n1632), .Z(n1186) );
  CND3X4 U1444 ( .A(n1188), .B(n1187), .C(n1186), .Z(n2274) );
  CNR2X4 U1445 ( .A(n2274), .B(\req_vec_rr[13][0] ), .Z(n1962) );
  CIVX2 U1446 ( .A(\req_vec_rr[13][2] ), .Z(n2376) );
  CNR2X1 U1447 ( .A(n2376), .B(\req_vec_rr[13][1] ), .Z(n1775) );
  CND2X1 U1448 ( .A(n1962), .B(n1775), .Z(n1203) );
  CAN2X1 U1449 ( .A(n2166), .B(n2403), .Z(n1191) );
  CIVX2 U1450 ( .A(n1189), .Z(n1190) );
  CND3X2 U1451 ( .A(n1192), .B(n1191), .C(n1190), .Z(n2277) );
  CND2X4 U1452 ( .A(n2276), .B(n2183), .Z(n1193) );
  CNR2X4 U1453 ( .A(n2277), .B(n1193), .Z(n1951) );
  CNR2X1 U1454 ( .A(n1072), .B(\req_vec_rr[14][1] ), .Z(n1781) );
  CND2X2 U1455 ( .A(n1951), .B(n1781), .Z(n1202) );
  CNR2X2 U1456 ( .A(n1197), .B(n1196), .Z(n1198) );
  CND2X4 U1457 ( .A(n1199), .B(n1198), .Z(n1526) );
  CNR2X1 U1458 ( .A(n2413), .B(n1524), .Z(n1200) );
  CND3X2 U1459 ( .A(n2144), .B(n1200), .C(n1526), .Z(n2273) );
  CIVX2 U1460 ( .A(\req_vec_rr[12][1] ), .Z(n2336) );
  CND2X1 U1461 ( .A(\req_vec_rr[12][2] ), .B(n2336), .Z(n1778) );
  CIVX2 U1462 ( .A(n1778), .Z(n1645) );
  CND2X1 U1463 ( .A(n1964), .B(n1645), .Z(n1201) );
  CND4X2 U1464 ( .A(n1204), .B(n1203), .C(n1201), .D(n1202), .Z(n1455) );
  CAN2X2 U1465 ( .A(\req_vec_rr[0][0] ), .B(\req_vec_rr[0][1] ), .Z(n1758) );
  CNR2IX2 U1466 ( .B(\req_vec_rr[0][0] ), .A(\req_vec_rr[0][1] ), .Z(n1717) );
  CANR2X1 U1467 ( .A(n1426), .B(n1758), .C(n1717), .D(n1428), .Z(n1206) );
  CNR2IX2 U1468 ( .B(\req_vec_rr[0][1] ), .A(\req_vec_rr[0][0] ), .Z(n1984) );
  CIVX2 U1469 ( .A(\req_vec_rr[0][0] ), .Z(n2323) );
  CIVX3 U1470 ( .A(\req_vec_rr[0][1] ), .Z(n2333) );
  CAN2X2 U1471 ( .A(n2323), .B(n2333), .Z(n1918) );
  CANR2X1 U1472 ( .A(n1384), .B(n1984), .C(n1918), .D(n1388), .Z(n1205) );
  CND3X2 U1473 ( .A(n1206), .B(n1205), .C(\req_vec_rr[0][2] ), .Z(n1210) );
  CANR2X1 U1474 ( .A(n1392), .B(n1984), .C(n1918), .D(n1393), .Z(n1207) );
  CIVX3 U1475 ( .A(\req_vec_rr[0][2] ), .Z(n2329) );
  CND3X2 U1476 ( .A(n1208), .B(n1207), .C(n2329), .Z(n1209) );
  CND3X4 U1477 ( .A(n1210), .B(n1209), .C(\req_vec_rr[0][3] ), .Z(n2297) );
  CANR2X1 U1478 ( .A(n1432), .B(n1984), .C(n1918), .D(n1341), .Z(n1212) );
  CANR2X1 U1479 ( .A(n1433), .B(n1717), .C(n1758), .D(n1434), .Z(n1211) );
  CND3X2 U1480 ( .A(n1212), .B(n1211), .C(\req_vec_rr[0][2] ), .Z(n1606) );
  CANR2X1 U1481 ( .A(n1441), .B(n1984), .C(n1918), .D(n1445), .Z(n1214) );
  CANR2X1 U1482 ( .A(n1440), .B(n1717), .C(n1758), .D(n1444), .Z(n1213) );
  CND3X2 U1483 ( .A(n1214), .B(n1213), .C(n2329), .Z(n1605) );
  CIVX1 U1484 ( .A(\req_vec_rr[0][3] ), .Z(n2299) );
  CND3X2 U1485 ( .A(n1606), .B(n1605), .C(n2299), .Z(n1215) );
  CND2X4 U1486 ( .A(n2297), .B(n1215), .Z(n2191) );
  CNIVX4 U1487 ( .A(n2191), .Z(n1695) );
  CND2X1 U1488 ( .A(\req_vec_rr[7][0] ), .B(\req_vec_rr[7][1] ), .Z(n1228) );
  CIVX2 U1489 ( .A(n1444), .Z(n1217) );
  CNR2X1 U1490 ( .A(\req_vec_rr[7][2] ), .B(\req_vec_rr[7][3] ), .Z(n1216) );
  COND1X1 U1491 ( .A(n1228), .B(n1217), .C(n1216), .Z(n1220) );
  CIVX3 U1492 ( .A(\req_vec_rr[7][1] ), .Z(n2340) );
  CIVX2 U1493 ( .A(\req_vec_rr[7][0] ), .Z(n1221) );
  CND2X1 U1494 ( .A(n2340), .B(n1221), .Z(n1230) );
  CNR2X1 U1495 ( .A(n1218), .B(n1230), .Z(n1219) );
  CNR2X1 U1496 ( .A(n1220), .B(n1219), .Z(n1225) );
  CNR2X2 U1497 ( .A(n1221), .B(\req_vec_rr[7][1] ), .Z(n1241) );
  CND2X1 U1498 ( .A(n1241), .B(n1365), .Z(n1224) );
  CNR2X2 U1499 ( .A(n2340), .B(\req_vec_rr[7][0] ), .Z(n1239) );
  CND2X1 U1500 ( .A(n1239), .B(n1222), .Z(n1223) );
  CND3X1 U1501 ( .A(n1225), .B(n1224), .C(n1223), .Z(n1235) );
  CIVX2 U1502 ( .A(n1241), .Z(n1245) );
  CIVX2 U1503 ( .A(n1239), .Z(n1247) );
  CNR2X1 U1504 ( .A(n1343), .B(n1247), .Z(n1226) );
  CNR2X1 U1505 ( .A(n1227), .B(n1226), .Z(n1233) );
  CIVX2 U1506 ( .A(n1228), .Z(n1251) );
  CIVX2 U1507 ( .A(\req_vec_rr[7][3] ), .Z(n2371) );
  CND2X1 U1508 ( .A(\req_vec_rr[7][2] ), .B(n2371), .Z(n1229) );
  CANR1X1 U1509 ( .A(n1373), .B(n1251), .C(n1229), .Z(n1232) );
  CIVX2 U1510 ( .A(n1230), .Z(n1252) );
  CND2X1 U1511 ( .A(n1252), .B(n1370), .Z(n1231) );
  CND3X2 U1512 ( .A(n1233), .B(n1232), .C(n1231), .Z(n1234) );
  CND2X2 U1513 ( .A(n1235), .B(n1234), .Z(n1259) );
  CND2X1 U1514 ( .A(n1393), .B(n1252), .Z(n1238) );
  CND2X1 U1515 ( .A(n1421), .B(n1251), .Z(n1237) );
  CNR2X1 U1516 ( .A(\req_vec_rr[7][2] ), .B(n2371), .Z(n1236) );
  CAN3X2 U1517 ( .A(n1238), .B(n1237), .C(n1236), .Z(n1244) );
  CND2X1 U1518 ( .A(n1239), .B(n1392), .Z(n1243) );
  CND2X1 U1519 ( .A(n1241), .B(n1240), .Z(n1242) );
  CND3X1 U1520 ( .A(n1244), .B(n1243), .C(n1242), .Z(n1257) );
  CNR2X1 U1521 ( .A(n1247), .B(n1246), .Z(n1248) );
  CNR2X1 U1522 ( .A(n1249), .B(n1248), .Z(n1255) );
  CNIVX2 U1523 ( .A(n1426), .Z(n1387) );
  CND2X1 U1524 ( .A(\req_vec_rr[7][2] ), .B(\req_vec_rr[7][3] ), .Z(n1250) );
  CANR1X1 U1525 ( .A(n1387), .B(n1251), .C(n1250), .Z(n1254) );
  CND2X1 U1526 ( .A(n1252), .B(n1427), .Z(n1253) );
  CND3X1 U1527 ( .A(n1255), .B(n1254), .C(n1253), .Z(n1256) );
  CND2X2 U1528 ( .A(n1257), .B(n1256), .Z(n1258) );
  CNR2X2 U1529 ( .A(n1259), .B(n1258), .Z(n1597) );
  CIVX2 U1530 ( .A(n1597), .Z(n2176) );
  CIVX3 U1531 ( .A(n2176), .Z(n2141) );
  CNR2X2 U1532 ( .A(n1695), .B(n2141), .Z(n1453) );
  CNR2IX1 U1533 ( .B(\req_vec_rr[4][1] ), .A(\req_vec_rr[4][0] ), .Z(n1286) );
  CND2X1 U1534 ( .A(n1392), .B(n1286), .Z(n1261) );
  CAN2X1 U1535 ( .A(\req_vec_rr[4][0] ), .B(\req_vec_rr[4][1] ), .Z(n1287) );
  CND2X1 U1536 ( .A(n1421), .B(n1287), .Z(n1260) );
  CND2X1 U1537 ( .A(n1261), .B(n1260), .Z(n1274) );
  CNR2X1 U1538 ( .A(\req_vec_rr[4][0] ), .B(\req_vec_rr[4][1] ), .Z(n1280) );
  CND2X1 U1539 ( .A(n1393), .B(n1280), .Z(n1264) );
  CNR2IX1 U1540 ( .B(\req_vec_rr[4][0] ), .A(\req_vec_rr[4][1] ), .Z(n1281) );
  CND2X1 U1541 ( .A(n1416), .B(n1281), .Z(n1263) );
  CIVX2 U1542 ( .A(\req_vec_rr[4][3] ), .Z(n2354) );
  CNR2X1 U1543 ( .A(\req_vec_rr[4][2] ), .B(n2354), .Z(n1262) );
  CND3X1 U1544 ( .A(n1264), .B(n1263), .C(n1262), .Z(n1273) );
  CND2X1 U1545 ( .A(n1425), .B(n1286), .Z(n1266) );
  CND2X2 U1546 ( .A(n1266), .B(n1265), .Z(n1267) );
  CIVX2 U1547 ( .A(n1267), .Z(n1271) );
  CND2X1 U1548 ( .A(\req_vec_rr[4][2] ), .B(\req_vec_rr[4][3] ), .Z(n1268) );
  CANR1X1 U1549 ( .A(n1281), .B(n1428), .C(n1268), .Z(n1270) );
  CND2X1 U1550 ( .A(n1388), .B(n1280), .Z(n1269) );
  CND3X2 U1551 ( .A(n1271), .B(n1270), .C(n1269), .Z(n1272) );
  COND1X2 U1552 ( .A(n1274), .B(n1273), .C(n1272), .Z(n1295) );
  CND2X1 U1553 ( .A(\req_vec_rr[4][2] ), .B(n2354), .Z(n1275) );
  CANR1X1 U1554 ( .A(n1281), .B(n1433), .C(n1275), .Z(n1279) );
  CND2X1 U1555 ( .A(n1435), .B(n1280), .Z(n1278) );
  CND2X1 U1556 ( .A(n1434), .B(n1287), .Z(n1277) );
  CND2X1 U1557 ( .A(n1432), .B(n1286), .Z(n1276) );
  CND4X2 U1558 ( .A(n1279), .B(n1278), .C(n1277), .D(n1276), .Z(n1293) );
  CND2X1 U1559 ( .A(n1445), .B(n1280), .Z(n1284) );
  CND2X2 U1560 ( .A(n1440), .B(n1281), .Z(n1283) );
  CNR2X1 U1561 ( .A(\req_vec_rr[4][2] ), .B(\req_vec_rr[4][3] ), .Z(n1282) );
  CND3X2 U1562 ( .A(n1284), .B(n1283), .C(n1282), .Z(n1285) );
  CIVX2 U1563 ( .A(n1285), .Z(n1291) );
  CND2X1 U1564 ( .A(n1441), .B(n1286), .Z(n1289) );
  CND2X2 U1565 ( .A(n1444), .B(n1287), .Z(n1288) );
  CAN2X1 U1566 ( .A(n1289), .B(n1288), .Z(n1290) );
  CND2X2 U1567 ( .A(n1291), .B(n1290), .Z(n1292) );
  CND2X2 U1568 ( .A(n1293), .B(n1292), .Z(n1294) );
  CNR2X4 U1569 ( .A(n1295), .B(n1294), .Z(n1466) );
  CIVX4 U1570 ( .A(\req_vec_rr[1][2] ), .Z(n2339) );
  CND2X2 U1571 ( .A(n2339), .B(\req_vec_rr[1][1] ), .Z(n1975) );
  CIVX4 U1572 ( .A(\req_vec_rr[1][1] ), .Z(n2374) );
  CND2X1 U1573 ( .A(n2374), .B(\req_vec_rr[1][2] ), .Z(n1798) );
  COND2X2 U1574 ( .A(n1296), .B(n1444), .C(n1433), .D(n1798), .Z(n1299) );
  CND2X1 U1575 ( .A(\req_vec_rr[1][1] ), .B(\req_vec_rr[1][2] ), .Z(n1927) );
  CIVX1 U1576 ( .A(\req_vec_rr[1][3] ), .Z(n2360) );
  CAN2X1 U1577 ( .A(\req_vec_rr[1][0] ), .B(n2360), .Z(n1297) );
  COND1X2 U1578 ( .A(n1434), .B(n1927), .C(n1297), .Z(n1298) );
  CNR2X4 U1579 ( .A(n1299), .B(n1298), .Z(n1302) );
  CIVX2 U1580 ( .A(n1440), .Z(n1300) );
  CND2X2 U1581 ( .A(n2374), .B(n2339), .Z(n1911) );
  CIVX2 U1582 ( .A(n1911), .Z(n2058) );
  CND2X1 U1583 ( .A(n1300), .B(n2058), .Z(n1301) );
  CND2X4 U1584 ( .A(n1302), .B(n1301), .Z(n1459) );
  CNR2X1 U1585 ( .A(\req_vec_rr[1][0] ), .B(\req_vec_rr[1][3] ), .Z(n1303) );
  CNR2X1 U1586 ( .A(n1432), .B(n1927), .Z(n1304) );
  CNR2X2 U1587 ( .A(n1305), .B(n1304), .Z(n1309) );
  CNR2X1 U1588 ( .A(n1445), .B(n1911), .Z(n1306) );
  CNR2X2 U1589 ( .A(n1307), .B(n1306), .Z(n1308) );
  CND2X2 U1590 ( .A(n1459), .B(n1460), .Z(n1546) );
  CNR2X4 U1591 ( .A(n1466), .B(n1546), .Z(n1355) );
  CNR3X1 U1592 ( .A(n1392), .B(\req_vec_rr[1][0] ), .C(n1975), .Z(n1312) );
  CIVDX1 U1593 ( .A(n1975), .Z0(n2115), .Z1(n1296) );
  CND2X1 U1594 ( .A(\req_vec_rr[1][0] ), .B(n2115), .Z(n1310) );
  CNR2X2 U1595 ( .A(n1312), .B(n1311), .Z(n1320) );
  CMXI2X1 U1596 ( .A0(n1393), .A1(n1416), .S(\req_vec_rr[1][0] ), .Z(n1313) );
  CND2X1 U1597 ( .A(n1313), .B(n2058), .Z(n1319) );
  CND3X1 U1598 ( .A(n1428), .B(\req_vec_rr[1][0] ), .C(n2374), .Z(n1317) );
  CNR2X1 U1599 ( .A(\req_vec_rr[1][0] ), .B(\req_vec_rr[1][1] ), .Z(n1315) );
  CND3X4 U1600 ( .A(n1318), .B(n1319), .C(n1320), .Z(n1660) );
  CIVX2 U1601 ( .A(\req_vec_rr[3][1] ), .Z(n2344) );
  CIVX2 U1602 ( .A(\req_vec_rr[3][0] ), .Z(n1322) );
  CNR2X2 U1603 ( .A(n2344), .B(n1322), .Z(n1345) );
  CND2X1 U1604 ( .A(n1345), .B(n1421), .Z(n1325) );
  CNR2X2 U1605 ( .A(n1322), .B(\req_vec_rr[3][1] ), .Z(n1346) );
  CANR1X1 U1606 ( .A(n1416), .B(n1346), .C(n1321), .Z(n1324) );
  CND2X1 U1607 ( .A(n1322), .B(\req_vec_rr[3][1] ), .Z(n1344) );
  CIVX2 U1608 ( .A(n1344), .Z(n1328) );
  CNR2X2 U1609 ( .A(\req_vec_rr[3][0] ), .B(\req_vec_rr[3][1] ), .Z(n1340) );
  CANR2X1 U1610 ( .A(n1392), .B(n1328), .C(n1340), .D(n1393), .Z(n1323) );
  CND3X2 U1611 ( .A(n1325), .B(n1324), .C(n1323), .Z(n1326) );
  CIVX3 U1612 ( .A(n1326), .Z(n1332) );
  CND2X1 U1613 ( .A(\req_vec_rr[3][2] ), .B(\req_vec_rr[3][3] ), .Z(n1327) );
  CANR1X1 U1614 ( .A(n1346), .B(n1428), .C(n1327), .Z(n1331) );
  CANR2X1 U1615 ( .A(n1426), .B(n1345), .C(n1328), .D(n1425), .Z(n1330) );
  CND2X1 U1616 ( .A(n1388), .B(n1340), .Z(n1329) );
  CNR2X4 U1617 ( .A(n1332), .B(n973), .Z(n1463) );
  CND2X1 U1618 ( .A(n1340), .B(n1445), .Z(n1333) );
  COND1X1 U1619 ( .A(n1344), .B(n1334), .C(n1333), .Z(n1339) );
  CND2X1 U1620 ( .A(n1345), .B(n1444), .Z(n1337) );
  CND2X1 U1621 ( .A(n1346), .B(n1440), .Z(n1336) );
  CNR2X1 U1622 ( .A(\req_vec_rr[3][2] ), .B(\req_vec_rr[3][3] ), .Z(n1335) );
  CND3X1 U1623 ( .A(n1337), .B(n1336), .C(n1335), .Z(n1338) );
  CNR2X2 U1624 ( .A(n1339), .B(n1338), .Z(n1353) );
  CND2X1 U1625 ( .A(n1341), .B(n1340), .Z(n1342) );
  CND2X1 U1626 ( .A(n1345), .B(n1434), .Z(n1349) );
  CND2X1 U1627 ( .A(n1346), .B(n1433), .Z(n1348) );
  CNR2IX1 U1628 ( .B(\req_vec_rr[3][2] ), .A(\req_vec_rr[3][3] ), .Z(n1347) );
  CND3X2 U1629 ( .A(n1349), .B(n1348), .C(n1347), .Z(n1350) );
  CNR2X2 U1630 ( .A(n1351), .B(n1350), .Z(n1352) );
  CNR2X4 U1631 ( .A(n1353), .B(n1352), .Z(n1464) );
  CND2X2 U1632 ( .A(n1463), .B(n1464), .Z(n1354) );
  CND3X4 U1633 ( .A(n1355), .B(n1660), .C(n1354), .Z(n1593) );
  CNR2IX1 U1634 ( .B(\req_vec_rr[6][0] ), .A(\req_vec_rr[6][1] ), .Z(n1374) );
  CIVX2 U1635 ( .A(\req_vec_rr[6][3] ), .Z(n2352) );
  CANR3X1 U1636 ( .A(n1374), .B(n1416), .C(\req_vec_rr[6][2] ), .D(n2352), .Z(
        n1359) );
  CIVX2 U1637 ( .A(\req_vec_rr[6][1] ), .Z(n1752) );
  CNR2X1 U1638 ( .A(n1752), .B(\req_vec_rr[6][0] ), .Z(n1376) );
  CND2X1 U1639 ( .A(n1376), .B(n1392), .Z(n1358) );
  CIVX2 U1640 ( .A(\req_vec_rr[6][0] ), .Z(n2334) );
  CNR2X2 U1641 ( .A(n1752), .B(n2334), .Z(n1372) );
  CND2X1 U1642 ( .A(n1372), .B(n1421), .Z(n1357) );
  CNR2X1 U1643 ( .A(\req_vec_rr[6][1] ), .B(\req_vec_rr[6][0] ), .Z(n1371) );
  CND2X1 U1644 ( .A(n1371), .B(n1420), .Z(n1356) );
  CND4X2 U1645 ( .A(n1359), .B(n1358), .C(n1357), .D(n1356), .Z(n1383) );
  CANR2X2 U1646 ( .A(n1361), .B(n1376), .C(n1360), .D(n1374), .Z(n1364) );
  CND2X1 U1647 ( .A(\req_vec_rr[6][2] ), .B(\req_vec_rr[6][3] ), .Z(n1362) );
  CANR1X2 U1648 ( .A(n1374), .B(n1365), .C(n975), .Z(n1369) );
  CANR3X1 U1649 ( .A(n1372), .B(n1444), .C(\req_vec_rr[6][3] ), .D(
        \req_vec_rr[6][2] ), .Z(n1368) );
  CND2X1 U1650 ( .A(n1371), .B(n1366), .Z(n1367) );
  CND3X2 U1651 ( .A(n1369), .B(n1368), .C(n1367), .Z(n1381) );
  CND2X1 U1652 ( .A(n1371), .B(n1370), .Z(n1379) );
  CANR2X2 U1653 ( .A(n1376), .B(n1375), .C(n1433), .D(n1374), .Z(n1377) );
  CND3X2 U1654 ( .A(n1379), .B(n1378), .C(n1377), .Z(n1380) );
  CND4X4 U1655 ( .A(n1383), .B(n1382), .C(n1381), .D(n1380), .Z(n1614) );
  CIVX2 U1656 ( .A(\req_vec_rr[5][0] ), .Z(n1385) );
  CNR2X1 U1657 ( .A(n1385), .B(\req_vec_rr[5][1] ), .Z(n1405) );
  CIVX2 U1658 ( .A(\req_vec_rr[5][1] ), .Z(n2372) );
  CNR2X1 U1659 ( .A(\req_vec_rr[5][0] ), .B(n2372), .Z(n1404) );
  CANR2X1 U1660 ( .A(n1405), .B(n1428), .C(n1404), .D(n1384), .Z(n1391) );
  CNR2X2 U1661 ( .A(n1385), .B(n2372), .Z(n1408) );
  CND2X1 U1662 ( .A(\req_vec_rr[5][2] ), .B(\req_vec_rr[5][3] ), .Z(n1386) );
  CNR2X2 U1663 ( .A(\req_vec_rr[5][0] ), .B(\req_vec_rr[5][1] ), .Z(n1406) );
  CND2X1 U1664 ( .A(n1406), .B(n1388), .Z(n1389) );
  CND3X2 U1665 ( .A(n1391), .B(n1390), .C(n1389), .Z(n1415) );
  CANR2X1 U1666 ( .A(n1416), .B(n1405), .C(n1392), .D(n1404), .Z(n1397) );
  CND2X1 U1667 ( .A(n1406), .B(n927), .Z(n1396) );
  CNR2X1 U1668 ( .A(\req_vec_rr[5][2] ), .B(n2319), .Z(n1395) );
  CND2X1 U1669 ( .A(n1408), .B(n1421), .Z(n1394) );
  CND4X2 U1670 ( .A(n1397), .B(n1396), .C(n1395), .D(n1394), .Z(n1414) );
  CIVX1 U1671 ( .A(\req_vec_rr[5][2] ), .Z(n1398) );
  CND2X1 U1672 ( .A(n2319), .B(n1398), .Z(n1399) );
  CANR1X2 U1673 ( .A(n1408), .B(n1400), .C(n1399), .Z(n1403) );
  CANR2X1 U1674 ( .A(n1405), .B(n1440), .C(n1441), .D(n1404), .Z(n1402) );
  CND2X1 U1675 ( .A(n1406), .B(n1445), .Z(n1401) );
  CND3X2 U1676 ( .A(n1403), .B(n1402), .C(n1401), .Z(n1413) );
  CANR2X1 U1677 ( .A(n1405), .B(n1433), .C(n1432), .D(n1404), .Z(n1411) );
  CND2X1 U1678 ( .A(n1406), .B(n1435), .Z(n1410) );
  CND2X1 U1679 ( .A(\req_vec_rr[5][2] ), .B(n2319), .Z(n1407) );
  CANR1X1 U1680 ( .A(n1434), .B(n1408), .C(n1407), .Z(n1409) );
  CND3X2 U1681 ( .A(n1411), .B(n1410), .C(n1409), .Z(n1412) );
  CND4X2 U1682 ( .A(n1415), .B(n1414), .C(n1413), .D(n1412), .Z(n1596) );
  CND2X2 U1683 ( .A(n1614), .B(n1596), .Z(n1470) );
  CIVX4 U1684 ( .A(\req_vec_rr[2][0] ), .Z(n2301) );
  CND2X1 U1685 ( .A(\req_vec_rr[2][1] ), .B(n2301), .Z(n1424) );
  CNR2X2 U1686 ( .A(\req_vec_rr[2][1] ), .B(n2301), .Z(n1439) );
  CIVX1 U1687 ( .A(n1439), .Z(n1417) );
  CND2IX1 U1688 ( .B(n1417), .A(n1416), .Z(n1418) );
  CNR2X2 U1689 ( .A(\req_vec_rr[2][1] ), .B(\req_vec_rr[2][0] ), .Z(n1446) );
  CND2X1 U1690 ( .A(n1446), .B(n1420), .Z(n1423) );
  CIVX2 U1691 ( .A(\req_vec_rr[2][1] ), .Z(n2193) );
  CNR2X2 U1692 ( .A(n2193), .B(n2301), .Z(n1443) );
  CND3X4 U1693 ( .A(n974), .B(n1423), .C(n1422), .Z(n1462) );
  CIVX2 U1694 ( .A(n1424), .Z(n1442) );
  CANR2X1 U1695 ( .A(n1426), .B(n1443), .C(n1442), .D(n1425), .Z(n1431) );
  CND2X1 U1696 ( .A(n1446), .B(n1427), .Z(n1430) );
  CIVX2 U1697 ( .A(\req_vec_rr[2][2] ), .Z(n2332) );
  CANR1X1 U1698 ( .A(n1439), .B(n1428), .C(n2332), .Z(n1429) );
  CND3X2 U1699 ( .A(n1431), .B(n1430), .C(n1429), .Z(n1461) );
  CND3X4 U1700 ( .A(n1462), .B(n1461), .C(n933), .Z(n1479) );
  CANR2X1 U1701 ( .A(n1439), .B(n1433), .C(n1442), .D(n1432), .Z(n1438) );
  CANR1X1 U1702 ( .A(n1434), .B(n1443), .C(n2332), .Z(n1437) );
  CND2X1 U1703 ( .A(n1446), .B(n1435), .Z(n1436) );
  CND3X1 U1704 ( .A(n1438), .B(n1437), .C(n1436), .Z(n1451) );
  CANR2X2 U1705 ( .A(n1441), .B(n1442), .C(n1440), .D(n1439), .Z(n1449) );
  CANR1X1 U1706 ( .A(n1444), .B(n1443), .C(\req_vec_rr[2][2] ), .Z(n1448) );
  CND2X1 U1707 ( .A(n1446), .B(n1445), .Z(n1447) );
  CND3X1 U1708 ( .A(n1449), .B(n1448), .C(n1447), .Z(n1450) );
  CIVX2 U1709 ( .A(n933), .Z(n1609) );
  CND3X2 U1710 ( .A(n1451), .B(n1450), .C(n1609), .Z(n1478) );
  CND2X4 U1711 ( .A(n1479), .B(n1478), .Z(n1592) );
  CNR2X2 U1712 ( .A(n1470), .B(n1592), .Z(n1452) );
  CND2IX2 U1713 ( .B(n1593), .A(n1452), .Z(n2142) );
  CIVX4 U1714 ( .A(n2142), .Z(n2177) );
  CND2X4 U1715 ( .A(n1453), .B(n2177), .Z(n1454) );
  CIVX16 U1716 ( .A(n1454), .Z(n2280) );
  COND1X2 U1717 ( .A(n1456), .B(n1455), .C(n2280), .Z(n1488) );
  CNR2X4 U1718 ( .A(n1593), .B(n1592), .Z(n1476) );
  CIVX4 U1719 ( .A(n1596), .Z(n1615) );
  CND2X2 U1720 ( .A(n1476), .B(n1615), .Z(n1457) );
  CIVX4 U1721 ( .A(n1457), .Z(n2283) );
  CNR2X1 U1722 ( .A(\req_vec_rr[5][0] ), .B(n2319), .Z(n1458) );
  CND2X2 U1723 ( .A(n2283), .B(n1458), .Z(n1981) );
  CND2X1 U1724 ( .A(\req_vec_rr[5][2] ), .B(n2372), .Z(n1796) );
  CIVX2 U1725 ( .A(n1796), .Z(n1654) );
  CND2X1 U1726 ( .A(n1972), .B(n1654), .Z(n1474) );
  CIVX4 U1727 ( .A(n1660), .Z(n2284) );
  CIVX2 U1728 ( .A(\req_vec_rr[1][0] ), .Z(n1659) );
  CND2X1 U1729 ( .A(n2284), .B(n1659), .Z(n1974) );
  CND2X4 U1730 ( .A(n1460), .B(n1459), .Z(n1607) );
  CND2X4 U1731 ( .A(n1480), .B(n1660), .Z(n2225) );
  CND3X2 U1732 ( .A(n1462), .B(n1461), .C(n934), .Z(n1656) );
  CNR2X2 U1733 ( .A(n2225), .B(n1656), .Z(n2285) );
  CND2X4 U1734 ( .A(n2285), .B(n2301), .Z(n1973) );
  CNR2X1 U1735 ( .A(\req_vec_rr[2][1] ), .B(n2332), .Z(n1799) );
  CIVX2 U1736 ( .A(n1799), .Z(n1550) );
  COND2X1 U1737 ( .A(n1798), .B(n1974), .C(n1973), .D(n1550), .Z(n1469) );
  CND2X4 U1738 ( .A(n1464), .B(n1463), .Z(n1465) );
  CIVX4 U1739 ( .A(n1465), .Z(n1602) );
  CNR2IX4 U1740 ( .B(n1466), .A(n1602), .Z(n2187) );
  CNR2X4 U1741 ( .A(n1592), .B(n2225), .Z(n2188) );
  CNR2X1 U1742 ( .A(n2354), .B(\req_vec_rr[4][0] ), .Z(n1467) );
  CND3X4 U1743 ( .A(n2187), .B(n2188), .C(n1467), .Z(n1977) );
  CIVX2 U1744 ( .A(\req_vec_rr[4][1] ), .Z(n2330) );
  CND2X1 U1745 ( .A(\req_vec_rr[4][2] ), .B(n2330), .Z(n1655) );
  CNR2X1 U1746 ( .A(n1977), .B(n1655), .Z(n1468) );
  COND1X2 U1747 ( .A(n1469), .B(n1468), .C(n1982), .Z(n1473) );
  CNR2X1 U1748 ( .A(\req_vec_rr[7][0] ), .B(n2371), .Z(n1905) );
  CNR2IX2 U1749 ( .B(n1597), .A(n1470), .Z(n1471) );
  CND2X4 U1750 ( .A(n1476), .B(n1471), .Z(n2291) );
  CNR2X1 U1751 ( .A(n2415), .B(\req_vec_rr[7][1] ), .Z(n1794) );
  COND3X1 U1752 ( .A(n1981), .B(n1474), .C(n1472), .D(n1473), .Z(n1486) );
  CNR2X2 U1753 ( .A(n1615), .B(n1614), .Z(n1475) );
  CND2X4 U1754 ( .A(n1476), .B(n1475), .Z(n2292) );
  CND2X1 U1755 ( .A(n2334), .B(\req_vec_rr[6][3] ), .Z(n1477) );
  CNR2X4 U1756 ( .A(n2292), .B(n1477), .Z(n1983) );
  CIVX2 U1757 ( .A(\req_vec_rr[6][2] ), .Z(n2400) );
  CNR2X1 U1758 ( .A(n2400), .B(\req_vec_rr[6][1] ), .Z(n1802) );
  CND3X1 U1759 ( .A(n1983), .B(n2293), .C(n1802), .Z(n1484) );
  CND2XL U1760 ( .A(n1922), .B(n1918), .Z(n1483) );
  CIVX2 U1761 ( .A(\req_vec_rr[3][3] ), .Z(n2348) );
  CNR2X1 U1762 ( .A(\req_vec_rr[3][0] ), .B(n2348), .Z(n1907) );
  CND2X4 U1763 ( .A(n1479), .B(n1478), .Z(n1548) );
  CND2X2 U1764 ( .A(n1480), .B(n1660), .Z(n1481) );
  CNR2X4 U1765 ( .A(n1548), .B(n1481), .Z(n1617) );
  CND2X4 U1766 ( .A(n1617), .B(n1602), .Z(n2282) );
  CNR2IX4 U1767 ( .B(n1907), .A(n2282), .Z(n1986) );
  CNR2X1 U1768 ( .A(\req_vec_rr[3][1] ), .B(n2232), .Z(n1801) );
  CND3XL U1769 ( .A(n1986), .B(n2293), .C(n1801), .Z(n1482) );
  CND3X1 U1770 ( .A(n1484), .B(n1483), .C(n1482), .Z(n1485) );
  CNR2X2 U1771 ( .A(n1486), .B(n1485), .Z(n1487) );
  CND2X2 U1772 ( .A(n1488), .B(n1487), .Z(gnt_nxt[12]) );
  CIVX2 U1773 ( .A(n2174), .Z(n1566) );
  CND2X4 U1774 ( .A(n1490), .B(n1489), .Z(n1570) );
  CNR2X4 U1775 ( .A(n1500), .B(n1570), .Z(n1498) );
  CND4X2 U1776 ( .A(n1494), .B(n1493), .C(n1492), .D(n1491), .Z(n1495) );
  CND2X2 U1777 ( .A(n1516), .B(n1495), .Z(n1496) );
  CIVX2 U1778 ( .A(n1496), .Z(n1497) );
  CNR3X2 U1779 ( .A(n938), .B(\req_vec_rr[15][0] ), .C(\req_vec_rr[15][3] ), 
        .Z(n1499) );
  CND2X2 U1780 ( .A(n1566), .B(n1499), .Z(n2080) );
  CNR2X1 U1781 ( .A(n2080), .B(n1774), .Z(n1538) );
  CIVX2 U1782 ( .A(n1642), .Z(n1777) );
  CNR2IX2 U1783 ( .B(n1516), .A(n1500), .Z(n1569) );
  CIVX4 U1784 ( .A(n2215), .Z(n2240) );
  CNR2X1 U1785 ( .A(\req_vec_rr[10][3] ), .B(\req_vec_rr[10][0] ), .Z(n1501)
         );
  CND2X4 U1786 ( .A(n2240), .B(n1501), .Z(n2084) );
  CND2X2 U1787 ( .A(n2082), .B(n1775), .Z(n1503) );
  COND1X1 U1788 ( .A(n1777), .B(n2084), .C(n1503), .Z(n1520) );
  CIVX2 U1789 ( .A(\req_vec_rr[8][1] ), .Z(n2335) );
  CND2X1 U1790 ( .A(n2335), .B(\req_vec_rr[8][2] ), .Z(n1784) );
  CND2X2 U1791 ( .A(n1505), .B(n1504), .Z(n1506) );
  CIVX2 U1792 ( .A(n1506), .Z(n1511) );
  CND2X2 U1793 ( .A(n1508), .B(n1507), .Z(n1509) );
  CIVX2 U1794 ( .A(n1509), .Z(n1510) );
  CND3X2 U1795 ( .A(n1511), .B(n1510), .C(\req_vec_rr[8][2] ), .Z(n1512) );
  CIVX2 U1796 ( .A(n1512), .Z(n1515) );
  CND2X1 U1797 ( .A(n1513), .B(n2328), .Z(n1514) );
  CND2IX2 U1798 ( .B(n1515), .A(n1514), .Z(n1582) );
  COND1X2 U1799 ( .A(\req_vec_rr[8][3] ), .B(n1582), .C(n1676), .Z(n2247) );
  CNR2X1 U1800 ( .A(\req_vec_rr[9][0] ), .B(\req_vec_rr[9][3] ), .Z(n1517) );
  CNR2IX2 U1801 ( .B(n1517), .A(n2268), .Z(n2087) );
  CND2X1 U1802 ( .A(n2087), .B(n1783), .Z(n1518) );
  COND1X1 U1803 ( .A(n1784), .B(n2089), .C(n1518), .Z(n1519) );
  CNR2X2 U1804 ( .A(n1520), .B(n1519), .Z(n1536) );
  CNR2XL U1805 ( .A(n2403), .B(\req_vec_rr[14][0] ), .Z(n1521) );
  CNR2IX2 U1806 ( .B(n1521), .A(n2175), .Z(n1523) );
  CNR2IX2 U1807 ( .B(n2166), .A(n1522), .Z(n2172) );
  CND2X2 U1808 ( .A(n1523), .B(n2172), .Z(n2094) );
  CND2IX1 U1809 ( .B(n2094), .A(n1781), .Z(n1535) );
  CNR2X1 U1810 ( .A(\req_vec_rr[12][3] ), .B(\req_vec_rr[12][0] ), .Z(n1527)
         );
  CIVX2 U1811 ( .A(n1524), .Z(n1525) );
  CND2X2 U1812 ( .A(n1526), .B(n1525), .Z(n1575) );
  CNR2IX2 U1813 ( .B(n1527), .A(n1575), .Z(n1528) );
  CND2X4 U1814 ( .A(n2276), .B(n1528), .Z(n2098) );
  CNR2X1 U1815 ( .A(n2098), .B(n1778), .Z(n1533) );
  CNR2X1 U1816 ( .A(n1529), .B(n1629), .Z(n1530) );
  CND2X2 U1817 ( .A(n1631), .B(n1530), .Z(n2212) );
  CNR2X1 U1818 ( .A(\req_vec_rr[11][0] ), .B(\req_vec_rr[11][3] ), .Z(n1531)
         );
  CND2X4 U1819 ( .A(n2271), .B(n1531), .Z(n2096) );
  CNR2X2 U1820 ( .A(n2096), .B(n1782), .Z(n1532) );
  CNR2X2 U1821 ( .A(n1533), .B(n1532), .Z(n1534) );
  CND3X2 U1822 ( .A(n1536), .B(n1535), .C(n1534), .Z(n1537) );
  COND1X2 U1823 ( .A(n1538), .B(n1537), .C(n2280), .Z(n1564) );
  CNR2X1 U1824 ( .A(\req_vec_rr[3][0] ), .B(\req_vec_rr[3][3] ), .Z(n2113) );
  CND2XL U1825 ( .A(n2113), .B(n1801), .Z(n1541) );
  CIVDX3 U1826 ( .A(n1607), .Z0(n1480), .Z1(n1539) );
  CND2X2 U1827 ( .A(n1539), .B(n1659), .Z(n2116) );
  CIVXL U1828 ( .A(n1798), .Z(n1661) );
  CND2IX1 U1829 ( .B(n2116), .A(n1661), .Z(n1540) );
  COND1X1 U1830 ( .A(n1541), .B(n2282), .C(n1540), .Z(n1543) );
  CNR2X1 U1831 ( .A(\req_vec_rr[0][3] ), .B(\req_vec_rr[0][0] ), .Z(n1542) );
  CND2X4 U1832 ( .A(n1838), .B(n1542), .Z(n2120) );
  CND2XL U1833 ( .A(n2333), .B(\req_vec_rr[0][2] ), .Z(n1797) );
  CNR2X1 U1834 ( .A(n2120), .B(n1797), .Z(n1558) );
  CNR2X2 U1835 ( .A(n1543), .B(n1558), .Z(n1555) );
  CNR2XL U1836 ( .A(\req_vec_rr[7][0] ), .B(\req_vec_rr[7][3] ), .Z(n1544) );
  CNR2IX4 U1837 ( .B(n1544), .A(n2291), .Z(n2112) );
  CND2X1 U1838 ( .A(n2112), .B(n1794), .Z(n1554) );
  CNR2X1 U1839 ( .A(\req_vec_rr[4][0] ), .B(\req_vec_rr[4][3] ), .Z(n1545) );
  CND3X2 U1840 ( .A(n2187), .B(n2188), .C(n1545), .Z(n2122) );
  CNR2X1 U1841 ( .A(n2122), .B(n1655), .Z(n1552) );
  CNR2X2 U1842 ( .A(n2284), .B(n1546), .Z(n1547) );
  CND2X4 U1843 ( .A(n1548), .B(n1547), .Z(n2228) );
  CIVX4 U1844 ( .A(n2228), .Z(n2147) );
  CNR2X1 U1845 ( .A(n934), .B(\req_vec_rr[2][0] ), .Z(n1549) );
  CND2X4 U1846 ( .A(n2147), .B(n1549), .Z(n2125) );
  CNR2X1 U1847 ( .A(n2125), .B(n1550), .Z(n1551) );
  CNR2X2 U1848 ( .A(n1552), .B(n1551), .Z(n1553) );
  CND3X2 U1849 ( .A(n1555), .B(n1554), .C(n1553), .Z(n1562) );
  CND2X1 U1850 ( .A(n2334), .B(n2352), .Z(n1556) );
  CNR2X4 U1851 ( .A(n2292), .B(n1556), .Z(n2107) );
  CND2X1 U1852 ( .A(n2107), .B(n1802), .Z(n1557) );
  CIVX2 U1853 ( .A(n1558), .Z(n1559) );
  CND2X1 U1854 ( .A(n1559), .B(n2236), .Z(n1560) );
  COND1X2 U1855 ( .A(n1562), .B(n1561), .C(n1560), .Z(n1563) );
  CND2X2 U1856 ( .A(n1564), .B(n1563), .Z(gnt_nxt[4]) );
  CNR3X2 U1857 ( .A(n938), .B(\req_vec_rr[15][3] ), .C(n2321), .Z(n1565) );
  CND2X2 U1858 ( .A(n1566), .B(n1565), .Z(n1863) );
  CND2X1 U1859 ( .A(n2317), .B(\req_vec_rr[15][1] ), .Z(n2079) );
  CNR2X1 U1860 ( .A(n1863), .B(n2079), .Z(n1591) );
  CIVX2 U1861 ( .A(n938), .Z(n1568) );
  CNR2X1 U1862 ( .A(n2403), .B(n2183), .Z(n1567) );
  CND3X2 U1863 ( .A(n1568), .B(n2172), .C(n1567), .Z(n1870) );
  CNR2X1 U1864 ( .A(n1743), .B(\req_vec_rr[14][2] ), .Z(n2093) );
  CND2IX1 U1865 ( .B(n1870), .A(n2093), .Z(n1589) );
  CND2X1 U1866 ( .A(\req_vec_rr[10][1] ), .B(n2262), .Z(n2085) );
  CIVX2 U1867 ( .A(n1569), .Z(n1572) );
  CND2X2 U1868 ( .A(n1570), .B(\req_vec_rr[10][0] ), .Z(n1571) );
  CNR2X4 U1869 ( .A(n1572), .B(n1571), .Z(n2160) );
  CND2X4 U1870 ( .A(n2160), .B(n2416), .Z(n1866) );
  CNR2IX4 U1871 ( .B(n1573), .A(n2175), .Z(n1864) );
  CNR2X1 U1872 ( .A(\req_vec_rr[13][2] ), .B(n2316), .Z(n2081) );
  CND2X2 U1873 ( .A(n1864), .B(n2081), .Z(n1574) );
  COND1X2 U1874 ( .A(n2085), .B(n1866), .C(n1574), .Z(n1578) );
  CIVX2 U1875 ( .A(n1575), .Z(n2143) );
  CIVX2 U1876 ( .A(\req_vec_rr[12][0] ), .Z(n2300) );
  CNR2X1 U1877 ( .A(\req_vec_rr[12][3] ), .B(n2300), .Z(n1576) );
  CND3X2 U1878 ( .A(n2144), .B(n2143), .C(n1576), .Z(n1867) );
  CNR2IX1 U1879 ( .B(\req_vec_rr[12][1] ), .A(\req_vec_rr[12][2] ), .Z(n1963)
         );
  CIVX1 U1880 ( .A(n1963), .Z(n2097) );
  CNR2X1 U1881 ( .A(n1867), .B(n2097), .Z(n1577) );
  CNR2X1 U1882 ( .A(n1635), .B(\req_vec_rr[11][3] ), .Z(n1579) );
  CND2X4 U1883 ( .A(n2271), .B(n1579), .Z(n1872) );
  CND2X1 U1884 ( .A(\req_vec_rr[11][1] ), .B(n1580), .Z(n2095) );
  CNR2X1 U1885 ( .A(n1872), .B(n2095), .Z(n1586) );
  CNR2IX1 U1886 ( .B(n2203), .A(\req_vec_rr[9][2] ), .Z(n2086) );
  CIVXL U1887 ( .A(n2086), .Z(n1584) );
  CNR2X2 U1888 ( .A(n2268), .B(n1628), .Z(n2161) );
  CND2X4 U1889 ( .A(n2161), .B(n2379), .Z(n1876) );
  CND2X1 U1890 ( .A(n2414), .B(n2314), .Z(n1581) );
  CNR2X2 U1891 ( .A(n1582), .B(n1581), .Z(n1874) );
  CND2X1 U1892 ( .A(n2328), .B(\req_vec_rr[8][1] ), .Z(n2090) );
  COND1X1 U1893 ( .A(n1584), .B(n1876), .C(n1583), .Z(n1585) );
  CNR2X2 U1894 ( .A(n1586), .B(n1585), .Z(n1587) );
  CND3X2 U1895 ( .A(n1589), .B(n1588), .C(n1587), .Z(n1590) );
  COND1X2 U1896 ( .A(n1591), .B(n1590), .C(n2280), .Z(n1626) );
  CNR2X1 U1897 ( .A(\req_vec_rr[5][2] ), .B(n2372), .Z(n1971) );
  CIVX2 U1898 ( .A(n1971), .Z(n2109) );
  CNR2X4 U1899 ( .A(n1593), .B(n1592), .Z(n1616) );
  CND2X2 U1900 ( .A(n1615), .B(\req_vec_rr[5][0] ), .Z(n1594) );
  CIVX2 U1901 ( .A(n1594), .Z(n1595) );
  CND2X2 U1902 ( .A(n1616), .B(n1595), .Z(n2152) );
  CND2X1 U1903 ( .A(n1614), .B(\req_vec_rr[7][0] ), .Z(n1598) );
  CNR2X2 U1904 ( .A(n1599), .B(n1598), .Z(n1600) );
  CND2X2 U1905 ( .A(n1600), .B(n1616), .Z(n2150) );
  CNR2X2 U1906 ( .A(n2150), .B(\req_vec_rr[7][3] ), .Z(n1825) );
  CNR2X1 U1907 ( .A(n2340), .B(\req_vec_rr[7][2] ), .Z(n2111) );
  CND2X1 U1908 ( .A(n2111), .B(n1825), .Z(n1601) );
  COND1X1 U1909 ( .A(n2109), .B(n1853), .C(n1601), .Z(n1624) );
  CNR2X1 U1910 ( .A(n2344), .B(\req_vec_rr[3][2] ), .Z(n2114) );
  CAN2X1 U1911 ( .A(n1602), .B(\req_vec_rr[3][0] ), .Z(n1603) );
  CND2X2 U1912 ( .A(n1603), .B(n1617), .Z(n2153) );
  CNR2IXL U1913 ( .B(\req_vec_rr[0][0] ), .A(\req_vec_rr[0][3] ), .Z(n1604) );
  CND3X1 U1914 ( .A(n1606), .B(n1605), .C(n1604), .Z(n1844) );
  CND2X1 U1915 ( .A(n2329), .B(\req_vec_rr[0][1] ), .Z(n2119) );
  CNR2X1 U1916 ( .A(n1844), .B(n2119), .Z(n1621) );
  CND2X2 U1917 ( .A(n1607), .B(\req_vec_rr[1][0] ), .Z(n1848) );
  CNR2XL U1918 ( .A(n1848), .B(n1975), .Z(n1608) );
  CNR2X2 U1919 ( .A(n1621), .B(n1608), .Z(n1612) );
  CND2X1 U1920 ( .A(\req_vec_rr[2][1] ), .B(n2332), .Z(n2124) );
  CND2X1 U1921 ( .A(n1609), .B(\req_vec_rr[2][0] ), .Z(n1827) );
  CNR2X1 U1922 ( .A(n2124), .B(n1827), .Z(n1610) );
  CANR1X2 U1923 ( .A(n2114), .B(n1831), .C(n1613), .Z(n1620) );
  CNR2X2 U1924 ( .A(n2151), .B(\req_vec_rr[6][3] ), .Z(n1832) );
  CNR2X1 U1925 ( .A(n1752), .B(\req_vec_rr[6][2] ), .Z(n2106) );
  CND2X1 U1926 ( .A(n1832), .B(n2106), .Z(n1619) );
  CND3X4 U1927 ( .A(n2187), .B(\req_vec_rr[4][0] ), .C(n1617), .Z(n2154) );
  CNR2X2 U1928 ( .A(n2154), .B(\req_vec_rr[4][3] ), .Z(n1854) );
  CNR2IX1 U1929 ( .B(\req_vec_rr[4][1] ), .A(\req_vec_rr[4][2] ), .Z(n1976) );
  CND2X1 U1930 ( .A(n1854), .B(n1976), .Z(n1618) );
  CND3X2 U1931 ( .A(n1620), .B(n1619), .C(n1618), .Z(n1623) );
  COND1X2 U1932 ( .A(n1624), .B(n1623), .C(n1622), .Z(n1625) );
  CND2X2 U1933 ( .A(n1626), .B(n1625), .Z(gnt_nxt[3]) );
  CND3X2 U1934 ( .A(n1627), .B(\req_vec_rr[15][0] ), .C(n2276), .Z(n1730) );
  CNR2X1 U1935 ( .A(n1730), .B(n1774), .Z(n1651) );
  CAN2X2 U1936 ( .A(n2160), .B(\req_vec_rr[10][3] ), .Z(n1708) );
  CNR2X2 U1937 ( .A(n1628), .B(n2379), .Z(n1736) );
  CIVX2 U1938 ( .A(n1629), .Z(n1630) );
  CND2X4 U1939 ( .A(n1631), .B(n1630), .Z(n1633) );
  CNR2X4 U1940 ( .A(n1633), .B(n1632), .Z(n1735) );
  CNR2X1 U1941 ( .A(n1635), .B(n1634), .Z(n1732) );
  CAN2XL U1942 ( .A(n1636), .B(n1732), .Z(n1637) );
  CND2X2 U1943 ( .A(n1735), .B(n1637), .Z(n1639) );
  CND3X2 U1944 ( .A(n1640), .B(n1639), .C(n1638), .Z(n1641) );
  CANR1X2 U1945 ( .A(n1642), .B(n1708), .C(n1641), .Z(n1649) );
  CND2IX1 U1946 ( .B(n1643), .A(\req_vec_rr[14][0] ), .Z(n1644) );
  CNR2X4 U1947 ( .A(n1644), .B(n2277), .Z(n1744) );
  CND2X1 U1948 ( .A(n1744), .B(n1781), .Z(n1648) );
  CNR2X4 U1949 ( .A(n2274), .B(n1889), .Z(n1745) );
  CND2X1 U1950 ( .A(n1745), .B(n1775), .Z(n1647) );
  CND2X1 U1951 ( .A(n1742), .B(n1645), .Z(n1646) );
  CND4X2 U1952 ( .A(n1649), .B(n1648), .C(n1647), .D(n1646), .Z(n1650) );
  COND1X2 U1953 ( .A(n1651), .B(n1650), .C(n2280), .Z(n1673) );
  CNR2X2 U1954 ( .A(n2151), .B(n2352), .Z(n1753) );
  CND2X1 U1955 ( .A(n1753), .B(n1802), .Z(n1653) );
  CNR2X2 U1956 ( .A(n2150), .B(n2371), .Z(n1762) );
  CND2X1 U1957 ( .A(n1762), .B(n1794), .Z(n1652) );
  CND2X2 U1958 ( .A(n1653), .B(n1652), .Z(n1671) );
  CNR2X4 U1959 ( .A(n2152), .B(n2319), .Z(n1755) );
  CND2X1 U1960 ( .A(n1755), .B(n1654), .Z(n1667) );
  CIVX2 U1961 ( .A(n1655), .Z(n1803) );
  CIVX2 U1962 ( .A(n1656), .Z(n1657) );
  CND2X2 U1963 ( .A(n1657), .B(\req_vec_rr[2][0] ), .Z(n1658) );
  CNR2X2 U1964 ( .A(n2225), .B(n1658), .Z(n1757) );
  CND2X1 U1965 ( .A(n1757), .B(n1799), .Z(n1663) );
  CND2X1 U1966 ( .A(n1922), .B(n1717), .Z(n1668) );
  CNR2X1 U1967 ( .A(n1660), .B(n1659), .Z(n1759) );
  CND2X1 U1968 ( .A(n1759), .B(n1661), .Z(n1662) );
  CND3X1 U1969 ( .A(n1663), .B(n1668), .C(n1662), .Z(n1664) );
  CANR1X1 U1970 ( .A(n1803), .B(n1754), .C(n1664), .Z(n1666) );
  CNR2X2 U1971 ( .A(n2153), .B(n2348), .Z(n1756) );
  CND2X1 U1972 ( .A(n1756), .B(n1801), .Z(n1665) );
  CND3X1 U1973 ( .A(n1667), .B(n1666), .C(n1665), .Z(n1670) );
  CND2X1 U1974 ( .A(n1668), .B(n2236), .Z(n1669) );
  COND1X2 U1975 ( .A(n1671), .B(n1670), .C(n1669), .Z(n1672) );
  CND2X2 U1976 ( .A(n1673), .B(n1672), .Z(gnt_nxt[13]) );
  CNR2X1 U1977 ( .A(n1730), .B(n2079), .Z(n1686) );
  CIVX2 U1978 ( .A(n2085), .Z(n1953) );
  CIVXL U1979 ( .A(n2095), .Z(n1674) );
  CAN2X1 U1980 ( .A(n1674), .B(n1732), .Z(n1675) );
  CND2X2 U1981 ( .A(n1735), .B(n1675), .Z(n1679) );
  CNIVX3 U1982 ( .A(n1676), .Z(n2267) );
  CNR2X2 U1983 ( .A(n2267), .B(\req_vec_rr[8][2] ), .Z(n1956) );
  CND2X1 U1984 ( .A(n1956), .B(n1731), .Z(n1678) );
  CND3X2 U1985 ( .A(n2204), .B(n2086), .C(n1736), .Z(n1677) );
  CND3X2 U1986 ( .A(n1679), .B(n1678), .C(n1677), .Z(n1680) );
  CANR1X2 U1987 ( .A(n1953), .B(n1708), .C(n1680), .Z(n1684) );
  CND2X1 U1988 ( .A(n1744), .B(n2093), .Z(n1683) );
  CND2X1 U1989 ( .A(n1742), .B(n1963), .Z(n1682) );
  CND2X1 U1990 ( .A(n1745), .B(n2081), .Z(n1681) );
  CND4X2 U1991 ( .A(n1684), .B(n1683), .C(n1682), .D(n1681), .Z(n1685) );
  COND1X2 U1992 ( .A(n1686), .B(n1685), .C(n2280), .Z(n1701) );
  CND2X1 U1993 ( .A(n1753), .B(n2106), .Z(n1688) );
  CND2X1 U1994 ( .A(n1762), .B(n2111), .Z(n1687) );
  CND2X2 U1995 ( .A(n1688), .B(n1687), .Z(n1699) );
  CNR2X1 U1996 ( .A(n2297), .B(\req_vec_rr[0][2] ), .Z(n1985) );
  CND2X1 U1997 ( .A(n1985), .B(n1758), .Z(n1696) );
  CND2X1 U1998 ( .A(n1759), .B(n2115), .Z(n1689) );
  CND3X2 U1999 ( .A(n1690), .B(n1696), .C(n1689), .Z(n1691) );
  CND2X1 U2000 ( .A(n1756), .B(n2114), .Z(n1692) );
  CND2X1 U2001 ( .A(n1696), .B(n2199), .Z(n1697) );
  COND1X2 U2002 ( .A(n1699), .B(n1698), .C(n1697), .Z(n1700) );
  CND2X2 U2003 ( .A(n1701), .B(n1700), .Z(gnt_nxt[11]) );
  CNR2X4 U2004 ( .A(gnt_nxt[13]), .B(gnt_nxt[11]), .Z(n1773) );
  CND2X1 U2005 ( .A(n2337), .B(n2317), .Z(n2038) );
  CNR2X1 U2006 ( .A(n1730), .B(n2038), .Z(n1714) );
  CNR2X1 U2007 ( .A(\req_vec_rr[10][1] ), .B(\req_vec_rr[10][2] ), .Z(n1891)
         );
  CNR2X1 U2008 ( .A(\req_vec_rr[11][1] ), .B(\req_vec_rr[11][2] ), .Z(n1871)
         );
  CAN2XL U2009 ( .A(n1732), .B(n1871), .Z(n1702) );
  CND2X2 U2010 ( .A(n1735), .B(n1702), .Z(n1706) );
  CND2X1 U2011 ( .A(n1956), .B(n1703), .Z(n1705) );
  CNR2X2 U2012 ( .A(n2203), .B(\req_vec_rr[9][2] ), .Z(n2042) );
  CND2X1 U2013 ( .A(n2204), .B(n979), .Z(n1704) );
  CND3X2 U2014 ( .A(n1704), .B(n1705), .C(n1706), .Z(n1707) );
  CANR1X2 U2015 ( .A(n1891), .B(n1708), .C(n1707), .Z(n1712) );
  CNR2X1 U2016 ( .A(\req_vec_rr[14][1] ), .B(\req_vec_rr[14][2] ), .Z(n2047)
         );
  CND2X1 U2017 ( .A(n1744), .B(n2047), .Z(n1711) );
  CNR2X1 U2018 ( .A(\req_vec_rr[13][2] ), .B(\req_vec_rr[13][1] ), .Z(n2039)
         );
  CND2X1 U2019 ( .A(n1745), .B(n2039), .Z(n1710) );
  CNR2X1 U2020 ( .A(\req_vec_rr[12][2] ), .B(\req_vec_rr[12][1] ), .Z(n1899)
         );
  CND2X1 U2021 ( .A(n1742), .B(n1899), .Z(n1709) );
  CND4X2 U2022 ( .A(n1712), .B(n1711), .C(n1710), .D(n1709), .Z(n1713) );
  COND1X2 U2023 ( .A(n1714), .B(n1713), .C(n2280), .Z(n1729) );
  CNR2X1 U2024 ( .A(\req_vec_rr[6][1] ), .B(\req_vec_rr[6][2] ), .Z(n2069) );
  CND2X1 U2025 ( .A(n1753), .B(n2069), .Z(n1716) );
  CNR2X1 U2026 ( .A(\req_vec_rr[7][1] ), .B(\req_vec_rr[7][2] ), .Z(n2061) );
  CND2X1 U2027 ( .A(n1762), .B(n2061), .Z(n1715) );
  CND2X2 U2028 ( .A(n1716), .B(n1715), .Z(n1727) );
  CNR2X1 U2029 ( .A(\req_vec_rr[5][2] ), .B(\req_vec_rr[5][1] ), .Z(n1845) );
  CND2X2 U2030 ( .A(n1755), .B(n1845), .Z(n1723) );
  CNR2X1 U2031 ( .A(\req_vec_rr[4][2] ), .B(\req_vec_rr[4][1] ), .Z(n1908) );
  CNR2X1 U2032 ( .A(\req_vec_rr[2][1] ), .B(\req_vec_rr[2][2] ), .Z(n1910) );
  CND2X1 U2033 ( .A(n1757), .B(n1910), .Z(n1719) );
  CND2X1 U2034 ( .A(n1985), .B(n1717), .Z(n1724) );
  CND2X1 U2035 ( .A(n1759), .B(n2058), .Z(n1718) );
  CND3X1 U2036 ( .A(n1719), .B(n1724), .C(n1718), .Z(n1720) );
  CANR1X1 U2037 ( .A(n1908), .B(n1754), .C(n1720), .Z(n1722) );
  CNR2X1 U2038 ( .A(\req_vec_rr[3][1] ), .B(\req_vec_rr[3][2] ), .Z(n2057) );
  CND2X1 U2039 ( .A(n1756), .B(n2057), .Z(n1721) );
  CND2X1 U2040 ( .A(n1724), .B(n2199), .Z(n1725) );
  COND1X2 U2041 ( .A(n1727), .B(n1726), .C(n1725), .Z(n1728) );
  CND2X2 U2042 ( .A(n1729), .B(n1728), .Z(gnt_nxt[9]) );
  CND2X1 U2043 ( .A(\req_vec_rr[15][1] ), .B(\req_vec_rr[15][2] ), .Z(n1995)
         );
  CNR2X1 U2044 ( .A(n1730), .B(n1995), .Z(n1751) );
  CND2X1 U2045 ( .A(\req_vec_rr[10][1] ), .B(\req_vec_rr[10][2] ), .Z(n1996)
         );
  CIVX2 U2046 ( .A(n1996), .Z(n1935) );
  CND3X1 U2047 ( .A(n2160), .B(\req_vec_rr[10][3] ), .C(n1935), .Z(n1740) );
  CND2X1 U2048 ( .A(\req_vec_rr[11][1] ), .B(\req_vec_rr[11][2] ), .Z(n2006)
         );
  CIVXL U2049 ( .A(n2006), .Z(n1733) );
  CAN2X1 U2050 ( .A(n1733), .B(n1732), .Z(n1734) );
  CND2X1 U2051 ( .A(n1735), .B(n1734), .Z(n1738) );
  CND2X1 U2052 ( .A(n2203), .B(\req_vec_rr[9][2] ), .Z(n1817) );
  CIVX2 U2053 ( .A(n1817), .Z(n2000) );
  CND3X1 U2054 ( .A(n2204), .B(n1736), .C(n2000), .Z(n1737) );
  CND4X1 U2055 ( .A(n1740), .B(n1739), .C(n1738), .D(n1737), .Z(n1741) );
  CIVX2 U2056 ( .A(n1741), .Z(n1749) );
  CND2X1 U2057 ( .A(\req_vec_rr[12][2] ), .B(\req_vec_rr[12][1] ), .Z(n2007)
         );
  CIVX2 U2058 ( .A(n2007), .Z(n1942) );
  CND2X1 U2059 ( .A(n1742), .B(n1942), .Z(n1748) );
  CNR2X1 U2060 ( .A(n1743), .B(n1072), .Z(n2005) );
  CND2X2 U2061 ( .A(n1744), .B(n2005), .Z(n1747) );
  CNR2X1 U2062 ( .A(n2376), .B(n2316), .Z(n1997) );
  CND2X1 U2063 ( .A(n1745), .B(n1997), .Z(n1746) );
  CND4X2 U2064 ( .A(n1749), .B(n1748), .C(n1747), .D(n1746), .Z(n1750) );
  COND1X2 U2065 ( .A(n1751), .B(n1750), .C(n2280), .Z(n1771) );
  CNR2X1 U2066 ( .A(n1752), .B(n2400), .Z(n2015) );
  CND2X1 U2067 ( .A(\req_vec_rr[5][2] ), .B(\req_vec_rr[5][1] ), .Z(n2017) );
  CIVX2 U2068 ( .A(n2017), .Z(n1926) );
  CND2X1 U2069 ( .A(\req_vec_rr[4][2] ), .B(\req_vec_rr[4][1] ), .Z(n2025) );
  CIVX2 U2070 ( .A(n2025), .Z(n1833) );
  CANR2X4 U2071 ( .A(n1755), .B(n1926), .C(n1833), .D(n1754), .Z(n1766) );
  CNR2X1 U2072 ( .A(n2344), .B(n2232), .Z(n2019) );
  CND2X1 U2073 ( .A(n1756), .B(n2019), .Z(n1765) );
  CND2X1 U2074 ( .A(\req_vec_rr[2][1] ), .B(\req_vec_rr[2][2] ), .Z(n2026) );
  CND2X1 U2075 ( .A(n1922), .B(n1758), .Z(n1767) );
  CIVXL U2076 ( .A(n1927), .Z(n2020) );
  CND2X1 U2077 ( .A(n1759), .B(n2020), .Z(n1760) );
  CAN3X2 U2078 ( .A(n1761), .B(n1767), .C(n1760), .Z(n1764) );
  CNR2X1 U2079 ( .A(n2340), .B(n2415), .Z(n2018) );
  CND4X2 U2080 ( .A(n1766), .B(n1765), .C(n1764), .D(n1763), .Z(n1769) );
  CND2X1 U2081 ( .A(n1767), .B(n2236), .Z(n1768) );
  COND1X2 U2082 ( .A(n976), .B(n1769), .C(n1768), .Z(n1770) );
  CND2X2 U2083 ( .A(n1771), .B(n1770), .Z(gnt_nxt[15]) );
  CNR2X4 U2084 ( .A(gnt_nxt[9]), .B(gnt_nxt[15]), .Z(n1772) );
  CND2X4 U2085 ( .A(n1772), .B(n1773), .Z(n2138) );
  CNR2X1 U2086 ( .A(n1863), .B(n1774), .Z(n1793) );
  CND2X2 U2087 ( .A(n1864), .B(n1775), .Z(n1776) );
  COND1X2 U2088 ( .A(n1777), .B(n1866), .C(n1776), .Z(n1780) );
  CNR2X1 U2089 ( .A(n1867), .B(n1778), .Z(n1779) );
  CNR2X2 U2090 ( .A(n1780), .B(n1779), .Z(n1791) );
  CND2IX1 U2091 ( .B(n1870), .A(n1781), .Z(n1790) );
  CNR2X1 U2092 ( .A(n1872), .B(n1782), .Z(n1788) );
  CIVXL U2093 ( .A(n1783), .Z(n1786) );
  COND1X1 U2094 ( .A(n1786), .B(n1876), .C(n1785), .Z(n1787) );
  CNR2X2 U2095 ( .A(n1788), .B(n1787), .Z(n1789) );
  CND3X2 U2096 ( .A(n1791), .B(n1790), .C(n1789), .Z(n1792) );
  COND1X2 U2097 ( .A(n1793), .B(n1792), .C(n2280), .Z(n1812) );
  CND2X1 U2098 ( .A(n1825), .B(n1794), .Z(n1795) );
  COND1X1 U2099 ( .A(n1796), .B(n1853), .C(n1795), .Z(n1810) );
  CNR2X1 U2100 ( .A(n1844), .B(n1797), .Z(n1807) );
  CNR2X2 U2101 ( .A(n2228), .B(n1827), .Z(n1850) );
  CND2X1 U2102 ( .A(n1832), .B(n1802), .Z(n1805) );
  CND2X1 U2103 ( .A(n1854), .B(n1803), .Z(n1804) );
  CND3X2 U2104 ( .A(n1806), .B(n1805), .C(n1804), .Z(n1809) );
  COND1X2 U2105 ( .A(n1810), .B(n1809), .C(n1808), .Z(n1811) );
  CND2X2 U2106 ( .A(n1812), .B(n1811), .Z(gnt_nxt[5]) );
  CNR2X1 U2107 ( .A(n1863), .B(n1995), .Z(n1824) );
  CND2X2 U2108 ( .A(n1864), .B(n1997), .Z(n1813) );
  COND1X2 U2109 ( .A(n1996), .B(n1866), .C(n1813), .Z(n1815) );
  CNR2X1 U2110 ( .A(n1867), .B(n2007), .Z(n1814) );
  CNR2X2 U2111 ( .A(n1815), .B(n1814), .Z(n1821) );
  CNR2X1 U2112 ( .A(n1872), .B(n2006), .Z(n1819) );
  CND2X1 U2113 ( .A(\req_vec_rr[8][1] ), .B(\req_vec_rr[8][2] ), .Z(n2002) );
  COND1X1 U2114 ( .A(n1817), .B(n1876), .C(n1816), .Z(n1818) );
  CNR2X2 U2115 ( .A(n1819), .B(n1818), .Z(n1820) );
  CND3X2 U2116 ( .A(n1822), .B(n1821), .C(n1820), .Z(n1823) );
  COND1X2 U2117 ( .A(n1824), .B(n1823), .C(n2280), .Z(n1843) );
  CNR2X1 U2118 ( .A(n1848), .B(n1927), .Z(n1826) );
  CND2XL U2119 ( .A(\req_vec_rr[0][1] ), .B(\req_vec_rr[0][2] ), .Z(n2023) );
  CNR2X2 U2120 ( .A(n1826), .B(n1837), .Z(n1829) );
  CND2X1 U2121 ( .A(n1829), .B(n1828), .Z(n1830) );
  CANR1X2 U2122 ( .A(n2019), .B(n1831), .C(n1830), .Z(n1836) );
  CND2X1 U2123 ( .A(n1832), .B(n2015), .Z(n1835) );
  CND2X1 U2124 ( .A(n1854), .B(n1833), .Z(n1834) );
  CND3X2 U2125 ( .A(n1836), .B(n1835), .C(n1834), .Z(n1840) );
  COND1X2 U2126 ( .A(n1841), .B(n1840), .C(n1839), .Z(n1842) );
  CND2X2 U2127 ( .A(n1843), .B(n1842), .Z(gnt_nxt[7]) );
  CNR2X4 U2128 ( .A(gnt_nxt[5]), .B(gnt_nxt[7]), .Z(n1888) );
  CND2X1 U2129 ( .A(n2333), .B(n2329), .Z(n2059) );
  CNR2X1 U2130 ( .A(n1844), .B(n2059), .Z(n1862) );
  CIVX2 U2131 ( .A(n1845), .Z(n2071) );
  CND2X2 U2132 ( .A(n1847), .B(n1846), .Z(n1852) );
  CNR2X1 U2133 ( .A(n1848), .B(n1911), .Z(n1849) );
  CANR3X1 U2134 ( .A(n1850), .B(n1910), .C(n1862), .D(n1849), .Z(n1851) );
  COND3X1 U2135 ( .A(n1853), .B(n2071), .C(n1852), .D(n1851), .Z(n1861) );
  CND2X1 U2136 ( .A(n1854), .B(n1908), .Z(n1859) );
  CIVXL U2137 ( .A(n2061), .Z(n1855) );
  COR3X1 U2138 ( .A(\req_vec_rr[7][3] ), .B(n1855), .C(n2150), .Z(n1858) );
  CIVXL U2139 ( .A(n2153), .Z(n1856) );
  CND3X1 U2140 ( .A(n1856), .B(n2057), .C(n2348), .Z(n1857) );
  CND3X2 U2141 ( .A(n1859), .B(n1858), .C(n1857), .Z(n1860) );
  COND2X2 U2142 ( .A(n1972), .B(n1862), .C(n1861), .D(n1860), .Z(n1886) );
  CNR2X1 U2143 ( .A(n1863), .B(n2038), .Z(n1884) );
  CIVX2 U2144 ( .A(n1891), .Z(n2041) );
  CND2X2 U2145 ( .A(n1864), .B(n2039), .Z(n1865) );
  COND1X2 U2146 ( .A(n2041), .B(n1866), .C(n1865), .Z(n1869) );
  CIVX1 U2147 ( .A(n1899), .Z(n2049) );
  CNR2X1 U2148 ( .A(n1867), .B(n2049), .Z(n1868) );
  CNR2X2 U2149 ( .A(n1869), .B(n1868), .Z(n1882) );
  CIVX2 U2150 ( .A(n1871), .Z(n2048) );
  CIVXL U2151 ( .A(n2042), .Z(n1877) );
  CND2X1 U2152 ( .A(n2335), .B(n2328), .Z(n2044) );
  CIVX2 U2153 ( .A(n2044), .Z(n1873) );
  CND2X1 U2154 ( .A(n1874), .B(n1873), .Z(n1875) );
  COND1X1 U2155 ( .A(n1877), .B(n1876), .C(n1875), .Z(n1878) );
  CNR2X2 U2156 ( .A(n1879), .B(n1878), .Z(n1880) );
  CND3X2 U2157 ( .A(n1882), .B(n1881), .C(n1880), .Z(n1883) );
  COND1X2 U2158 ( .A(n1884), .B(n1883), .C(n2280), .Z(n1885) );
  CND2X2 U2159 ( .A(n1886), .B(n1885), .Z(gnt_nxt[1]) );
  CNR2X4 U2160 ( .A(gnt_nxt[1]), .B(gnt_nxt[3]), .Z(n1887) );
  CND2X4 U2161 ( .A(n1888), .B(n1887), .Z(n2137) );
  CNR2X4 U2162 ( .A(n2138), .B(n2137), .Z(n2266) );
  CND2XL U2163 ( .A(n2039), .B(n1889), .Z(n1890) );
  CND2X1 U2164 ( .A(n1956), .B(n1892), .Z(n1893) );
  CND3X2 U2165 ( .A(n1895), .B(n1894), .C(n1893), .Z(n1897) );
  CNR2X2 U2166 ( .A(n1952), .B(n2048), .Z(n1896) );
  CNR3X4 U2167 ( .A(n1898), .B(n1897), .C(n1896), .Z(n1902) );
  CND2X1 U2168 ( .A(n1951), .B(n2047), .Z(n1901) );
  CND2X1 U2169 ( .A(n1964), .B(n1899), .Z(n1900) );
  CND3X2 U2170 ( .A(n1902), .B(n1901), .C(n1900), .Z(n1903) );
  COND1X2 U2171 ( .A(n1904), .B(n1903), .C(n2280), .Z(n1921) );
  CND2XL U2172 ( .A(n2061), .B(n1905), .Z(n1906) );
  CNR2X1 U2173 ( .A(n2291), .B(n1906), .Z(n1914) );
  CND2X1 U2174 ( .A(n2057), .B(n1907), .Z(n1909) );
  CIVX1 U2175 ( .A(n1908), .Z(n2062) );
  COND2X2 U2176 ( .A(n1909), .B(n2282), .C(n1977), .D(n2062), .Z(n1913) );
  CIVX2 U2177 ( .A(n1910), .Z(n2063) );
  COND2X1 U2178 ( .A(n1911), .B(n1974), .C(n1973), .D(n2063), .Z(n1912) );
  CNR3X2 U2179 ( .A(n1914), .B(n1913), .C(n1912), .Z(n1916) );
  CND2X1 U2180 ( .A(n1983), .B(n2069), .Z(n1915) );
  COND3X1 U2181 ( .A(n1981), .B(n2071), .C(n1916), .D(n1915), .Z(n1917) );
  CND2X2 U2182 ( .A(n1917), .B(n2293), .Z(n1920) );
  CND2X1 U2183 ( .A(n1985), .B(n1918), .Z(n1919) );
  CND3X2 U2184 ( .A(n1921), .B(n1920), .C(n1919), .Z(gnt_nxt[8]) );
  CND3X1 U2185 ( .A(n1983), .B(n1972), .C(n2015), .Z(n1925) );
  CND2XL U2186 ( .A(n1922), .B(n1984), .Z(n1924) );
  CND3XL U2187 ( .A(n1986), .B(n1972), .C(n2019), .Z(n1923) );
  CND3X1 U2188 ( .A(n1925), .B(n1924), .C(n1923), .Z(n1934) );
  CND2X1 U2189 ( .A(n1972), .B(n1926), .Z(n1932) );
  COND2X1 U2190 ( .A(n1927), .B(n1974), .C(n1973), .D(n2026), .Z(n1929) );
  CNR2X1 U2191 ( .A(n1977), .B(n2025), .Z(n1928) );
  COND1X2 U2192 ( .A(n1929), .B(n1928), .C(n1972), .Z(n1930) );
  COND3X1 U2193 ( .A(n1981), .B(n1932), .C(n1931), .D(n1930), .Z(n1933) );
  CNR2X2 U2194 ( .A(n1934), .B(n1933), .Z(n1950) );
  CND2X1 U2195 ( .A(n1962), .B(n1997), .Z(n1945) );
  CNR2X1 U2196 ( .A(n2006), .B(n1952), .Z(n1941) );
  CND3X1 U2197 ( .A(n2270), .B(n1935), .C(n2322), .Z(n1939) );
  CND2X1 U2198 ( .A(n1936), .B(n1955), .Z(n1937) );
  CND3X2 U2199 ( .A(n1939), .B(n1938), .C(n1937), .Z(n1940) );
  CNR2X2 U2200 ( .A(n1941), .B(n1940), .Z(n1944) );
  CND2X1 U2201 ( .A(n1964), .B(n1942), .Z(n1943) );
  CND4X2 U2202 ( .A(n1946), .B(n1944), .C(n1945), .D(n1943), .Z(n1947) );
  COND1X2 U2203 ( .A(n1948), .B(n1947), .C(n2280), .Z(n1949) );
  CND2X2 U2204 ( .A(n1950), .B(n1949), .Z(gnt_nxt[14]) );
  CNR2X4 U2205 ( .A(gnt_nxt[14]), .B(gnt_nxt[12]), .Z(n1993) );
  CND2X1 U2206 ( .A(n1951), .B(n2093), .Z(n1968) );
  CNR2X1 U2207 ( .A(n1952), .B(n2095), .Z(n1961) );
  CND3X1 U2208 ( .A(n2270), .B(n1953), .C(n2322), .Z(n1959) );
  CND3X1 U2209 ( .A(n2204), .B(n2086), .C(n1954), .Z(n1958) );
  CND2X1 U2210 ( .A(n1956), .B(n1955), .Z(n1957) );
  CND3X1 U2211 ( .A(n1959), .B(n1958), .C(n1957), .Z(n1960) );
  CNR2X2 U2212 ( .A(n1961), .B(n1960), .Z(n1967) );
  CND2X1 U2213 ( .A(n1962), .B(n2081), .Z(n1966) );
  CND2X1 U2214 ( .A(n1964), .B(n1963), .Z(n1965) );
  COND1X2 U2215 ( .A(n1970), .B(n1969), .C(n2280), .Z(n1991) );
  COND2X1 U2216 ( .A(n1975), .B(n1974), .C(n1973), .D(n2124), .Z(n1979) );
  CIVX1 U2217 ( .A(n1976), .Z(n2123) );
  CNR2X1 U2218 ( .A(n1977), .B(n2123), .Z(n1978) );
  CND3X1 U2219 ( .A(n1983), .B(n1982), .C(n2106), .Z(n1987) );
  CNR2X2 U2220 ( .A(n1989), .B(n1988), .Z(n1990) );
  CND2X2 U2221 ( .A(n1991), .B(n1990), .Z(gnt_nxt[10]) );
  CIVX3 U2222 ( .A(gnt_nxt[10]), .Z(n1992) );
  CND3X4 U2223 ( .A(n1994), .B(n1993), .C(n1992), .Z(n2140) );
  CNR2X1 U2224 ( .A(n1995), .B(n2080), .Z(n2014) );
  CND2X1 U2225 ( .A(n2082), .B(n1997), .Z(n1998) );
  CND2X2 U2226 ( .A(n1999), .B(n1998), .Z(n2004) );
  CND2X1 U2227 ( .A(n2087), .B(n2000), .Z(n2001) );
  COND1X1 U2228 ( .A(n2089), .B(n2002), .C(n2001), .Z(n2003) );
  CNR2X4 U2229 ( .A(n2004), .B(n2003), .Z(n2012) );
  CND2IX1 U2230 ( .B(n2094), .A(n2005), .Z(n2011) );
  CNR2X1 U2231 ( .A(n2096), .B(n2006), .Z(n2009) );
  CNR2X1 U2232 ( .A(n2098), .B(n2007), .Z(n2008) );
  CNR2X2 U2233 ( .A(n2009), .B(n2008), .Z(n2010) );
  CND3X2 U2234 ( .A(n2012), .B(n2011), .C(n2010), .Z(n2013) );
  COND1X2 U2235 ( .A(n2014), .B(n2013), .C(n2280), .Z(n2037) );
  CND2X1 U2236 ( .A(n2107), .B(n2015), .Z(n2016) );
  COND1X2 U2237 ( .A(n2110), .B(n2017), .C(n2016), .Z(n2035) );
  CND2X1 U2238 ( .A(n2112), .B(n2018), .Z(n2031) );
  CND2XL U2239 ( .A(n2019), .B(n2113), .Z(n2022) );
  CND2IX1 U2240 ( .B(n2116), .A(n2020), .Z(n2021) );
  COND1X1 U2241 ( .A(n2022), .B(n2282), .C(n2021), .Z(n2024) );
  CNR2X1 U2242 ( .A(n2120), .B(n2023), .Z(n2032) );
  CNR2X1 U2243 ( .A(n2024), .B(n2032), .Z(n2030) );
  CNR2X1 U2244 ( .A(n2025), .B(n2122), .Z(n2028) );
  CNR2X1 U2245 ( .A(n2125), .B(n2026), .Z(n2027) );
  CNR2X1 U2246 ( .A(n2028), .B(n2027), .Z(n2029) );
  COND1X2 U2247 ( .A(n2035), .B(n2034), .C(n2033), .Z(n2036) );
  CNR2X4 U2248 ( .A(gnt_nxt[6]), .B(gnt_nxt[4]), .Z(n2136) );
  CNR2X1 U2249 ( .A(n2038), .B(n2080), .Z(n2056) );
  CND2X2 U2250 ( .A(n2082), .B(n2039), .Z(n2040) );
  COND1X2 U2251 ( .A(n2041), .B(n2084), .C(n2040), .Z(n2046) );
  CND2X1 U2252 ( .A(n2087), .B(n2042), .Z(n2043) );
  COND1X1 U2253 ( .A(n2044), .B(n2089), .C(n2043), .Z(n2045) );
  CND2IX1 U2254 ( .B(n2094), .A(n2047), .Z(n2053) );
  CNR2X1 U2255 ( .A(n2096), .B(n2048), .Z(n2051) );
  CNR2X1 U2256 ( .A(n2098), .B(n2049), .Z(n2050) );
  CNR2X2 U2257 ( .A(n2051), .B(n2050), .Z(n2052) );
  CND3X2 U2258 ( .A(n2054), .B(n2053), .C(n2052), .Z(n2055) );
  COND1X2 U2259 ( .A(n2056), .B(n2055), .C(n2280), .Z(n2078) );
  CNR2X1 U2260 ( .A(n2120), .B(n2059), .Z(n2072) );
  CND2X1 U2261 ( .A(n2112), .B(n2061), .Z(n2067) );
  CNR2X1 U2262 ( .A(n2122), .B(n2062), .Z(n2065) );
  CNR2X1 U2263 ( .A(n2125), .B(n2063), .Z(n2064) );
  CNR2X1 U2264 ( .A(n2065), .B(n2064), .Z(n2066) );
  CND2X1 U2265 ( .A(n2107), .B(n2069), .Z(n2070) );
  COND1X1 U2266 ( .A(n2071), .B(n2110), .C(n2070), .Z(n2075) );
  CIVX2 U2267 ( .A(n2072), .Z(n2073) );
  CND2X1 U2268 ( .A(n2073), .B(n2236), .Z(n2074) );
  COND1X2 U2269 ( .A(n2076), .B(n2075), .C(n2074), .Z(n2077) );
  CND2X2 U2270 ( .A(n2078), .B(n2077), .Z(gnt_nxt[0]) );
  CNR2X1 U2271 ( .A(n2080), .B(n2079), .Z(n2105) );
  CND2X2 U2272 ( .A(n2082), .B(n2081), .Z(n2083) );
  CND2X1 U2273 ( .A(n2087), .B(n2086), .Z(n2088) );
  COND1X1 U2274 ( .A(n2090), .B(n2089), .C(n2088), .Z(n2091) );
  CNR2X2 U2275 ( .A(n2092), .B(n2091), .Z(n2103) );
  CND2IX1 U2276 ( .B(n2094), .A(n2093), .Z(n2102) );
  CNR2X1 U2277 ( .A(n2096), .B(n2095), .Z(n2100) );
  CNR2X1 U2278 ( .A(n2098), .B(n2097), .Z(n2099) );
  CNR2X2 U2279 ( .A(n2100), .B(n2099), .Z(n2101) );
  CND3X2 U2280 ( .A(n2103), .B(n2102), .C(n2101), .Z(n2104) );
  COND1X2 U2281 ( .A(n2105), .B(n2104), .C(n2280), .Z(n2134) );
  CND2X2 U2282 ( .A(n2107), .B(n2106), .Z(n2108) );
  COND1X2 U2283 ( .A(n2110), .B(n2109), .C(n2108), .Z(n2132) );
  CND2XL U2284 ( .A(n2114), .B(n2113), .Z(n2118) );
  CND2IX1 U2285 ( .B(n2116), .A(n2115), .Z(n2117) );
  COND1X1 U2286 ( .A(n2118), .B(n2282), .C(n2117), .Z(n2121) );
  CNR2X1 U2287 ( .A(n2120), .B(n2119), .Z(n2129) );
  CNR2X1 U2288 ( .A(n2123), .B(n2122), .Z(n2127) );
  CNR2X1 U2289 ( .A(n2125), .B(n2124), .Z(n2126) );
  CNR2X1 U2290 ( .A(n2127), .B(n2126), .Z(n2128) );
  COND1X2 U2291 ( .A(n2132), .B(n2131), .C(n2130), .Z(n2133) );
  CND2X2 U2292 ( .A(n2134), .B(n2133), .Z(gnt_nxt[2]) );
  CNR2X4 U2293 ( .A(gnt_nxt[0]), .B(gnt_nxt[2]), .Z(n2135) );
  CND2X4 U2294 ( .A(n2136), .B(n2135), .Z(n2139) );
  CNR2X4 U2295 ( .A(n2140), .B(n2139), .Z(n2265) );
  CND2X4 U2296 ( .A(n2266), .B(n2265), .Z(n2398) );
  CNR2X4 U2297 ( .A(n2138), .B(n2137), .Z(n2264) );
  CNR2X4 U2298 ( .A(n2140), .B(n2139), .Z(n2263) );
  CND2X4 U2299 ( .A(n2264), .B(n2263), .Z(n2303) );
  CNR2X2 U2300 ( .A(n2142), .B(n2141), .Z(n2167) );
  CND2X2 U2301 ( .A(n2144), .B(n2143), .Z(n2244) );
  CIVXL U2302 ( .A(n2244), .Z(n2145) );
  CND3X1 U2303 ( .A(n2167), .B(\req_vec_rr[12][0] ), .C(n2145), .Z(n2159) );
  CND2X1 U2304 ( .A(n2147), .B(\req_vec_rr[2][0] ), .Z(n2148) );
  CAN3X2 U2305 ( .A(n2150), .B(n2149), .C(n2148), .Z(n2158) );
  CND2X1 U2306 ( .A(n2152), .B(n2151), .Z(n2156) );
  CNR2X2 U2307 ( .A(n2156), .B(n2155), .Z(n2157) );
  CNR2X1 U2308 ( .A(n2161), .B(n2160), .Z(n2164) );
  CND2X1 U2309 ( .A(n2271), .B(\req_vec_rr[11][0] ), .Z(n2163) );
  CND2XL U2310 ( .A(n2247), .B(n2314), .Z(n2162) );
  CND3X2 U2311 ( .A(n2165), .B(n2177), .C(n2176), .Z(n2169) );
  CNR2X2 U2312 ( .A(n938), .B(n2166), .Z(n2250) );
  CND3X1 U2313 ( .A(n2167), .B(\req_vec_rr[13][0] ), .C(n2250), .Z(n2168) );
  CND2X2 U2314 ( .A(n2169), .B(n2168), .Z(n2170) );
  CIVX2 U2315 ( .A(n2172), .Z(n2173) );
  CNR2X2 U2316 ( .A(n938), .B(n2173), .Z(n2252) );
  CND4X1 U2317 ( .A(n2252), .B(n2177), .C(\req_vec_rr[14][0] ), .D(n2176), .Z(
        n2179) );
  CNR2X2 U2318 ( .A(n938), .B(n2174), .Z(n2251) );
  CND4X1 U2319 ( .A(n2177), .B(n2251), .C(\req_vec_rr[15][0] ), .D(n2176), .Z(
        n2178) );
  CND3X4 U2320 ( .A(n2180), .B(n2179), .C(n2178), .Z(n2182) );
  CND2X4 U2321 ( .A(n2182), .B(n2181), .Z(n2326) );
  CND2X4 U2322 ( .A(n2303), .B(n2320), .Z(n2369) );
  COND1XL U2323 ( .A(n2183), .B(n2398), .C(n2369), .Z(\req_vec_rr_d[14][0] )
         );
  CND2X2 U2324 ( .A(n2184), .B(\req_vec_rr[6][1] ), .Z(n2186) );
  CND2X2 U2325 ( .A(n2283), .B(\req_vec_rr[5][1] ), .Z(n2185) );
  CND2X2 U2326 ( .A(n2186), .B(n2185), .Z(n2202) );
  CNIVX4 U2327 ( .A(n2187), .Z(n2189) );
  CND2X4 U2328 ( .A(n2189), .B(n2188), .Z(n2190) );
  CIVX4 U2329 ( .A(n2190), .Z(n2286) );
  CIVDX1 U2330 ( .A(n2191), .Z0(n2227), .Z1(n1838) );
  CND2X1 U2331 ( .A(n2225), .B(\req_vec_rr[1][1] ), .Z(n2192) );
  COND3X1 U2332 ( .A(n2193), .B(n2228), .C(n2227), .D(n2192), .Z(n2194) );
  CANR1X2 U2333 ( .A(\req_vec_rr[4][1] ), .B(n2286), .C(n2194), .Z(n2198) );
  CNR2IX2 U2334 ( .B(\req_vec_rr[7][1] ), .A(n2291), .Z(n2196) );
  CNR2IX2 U2335 ( .B(\req_vec_rr[3][1] ), .A(n2282), .Z(n2195) );
  CNR2X2 U2336 ( .A(n2196), .B(n2195), .Z(n2197) );
  CND2X2 U2337 ( .A(n2199), .B(n2333), .Z(n2200) );
  COND1X4 U2338 ( .A(n2202), .B(n2201), .C(n2200), .Z(n2223) );
  CND2X1 U2339 ( .A(n2251), .B(\req_vec_rr[15][1] ), .Z(n2210) );
  CND2X1 U2340 ( .A(n2252), .B(\req_vec_rr[14][1] ), .Z(n2209) );
  CND2X1 U2341 ( .A(n2247), .B(\req_vec_rr[8][1] ), .Z(n2206) );
  CND2X1 U2342 ( .A(n2204), .B(n2203), .Z(n2205) );
  CND2X1 U2343 ( .A(n2206), .B(n2205), .Z(n2207) );
  CANR1X2 U2344 ( .A(\req_vec_rr[13][1] ), .B(n2250), .C(n2207), .Z(n2208) );
  CND3X2 U2345 ( .A(n2210), .B(n2209), .C(n2208), .Z(n2211) );
  CIVDX4 U2346 ( .A(n2212), .Z0(n2271), .Z1(n2213) );
  CNR2X4 U2347 ( .A(n2213), .B(n2342), .Z(n2214) );
  CIVX3 U2348 ( .A(n2214), .Z(n2219) );
  COR2X1 U2349 ( .A(n2244), .B(n2336), .Z(n2218) );
  COR2X1 U2350 ( .A(n2216), .B(n2215), .Z(n2217) );
  CND3X4 U2351 ( .A(n2219), .B(n2218), .C(n2217), .Z(n2220) );
  CND2X4 U2352 ( .A(n2220), .B(n2280), .Z(n2221) );
  CND3X4 U2353 ( .A(n2223), .B(n2222), .C(n2221), .Z(n2260) );
  CNR2X4 U2354 ( .A(n2224), .B(n2326), .Z(n2389) );
  COR2X1 U2355 ( .A(n2400), .B(n2292), .Z(n2231) );
  COND3X1 U2356 ( .A(n2228), .B(n2332), .C(n2227), .D(n2226), .Z(n2229) );
  CND2X2 U2357 ( .A(n2231), .B(n2230), .Z(n2239) );
  CND2X1 U2358 ( .A(n2283), .B(\req_vec_rr[5][2] ), .Z(n2235) );
  COND2X2 U2359 ( .A(n2232), .B(n2282), .C(n2291), .D(n2415), .Z(n2233) );
  CIVX2 U2360 ( .A(n2233), .Z(n2234) );
  CND2X2 U2361 ( .A(n2235), .B(n2234), .Z(n2238) );
  CND2X1 U2362 ( .A(n2236), .B(n2329), .Z(n2237) );
  CND2X1 U2363 ( .A(n2271), .B(\req_vec_rr[11][2] ), .Z(n2242) );
  CND2X1 U2364 ( .A(n2240), .B(\req_vec_rr[10][2] ), .Z(n2241) );
  CND2X2 U2365 ( .A(n2242), .B(n2241), .Z(n2246) );
  CNR2X1 U2366 ( .A(n2244), .B(n2243), .Z(n2245) );
  CNR2X2 U2367 ( .A(n2246), .B(n2245), .Z(n2256) );
  CND2XL U2368 ( .A(n2247), .B(\req_vec_rr[8][2] ), .Z(n2248) );
  COND1XL U2369 ( .A(n2357), .B(n2268), .C(n2248), .Z(n2249) );
  CANR1X1 U2370 ( .A(\req_vec_rr[13][2] ), .B(n2250), .C(n2249), .Z(n2255) );
  CND2X1 U2371 ( .A(n2251), .B(\req_vec_rr[15][2] ), .Z(n2254) );
  CND4X2 U2372 ( .A(n2256), .B(n2255), .C(n2254), .D(n2253), .Z(n2257) );
  CND2X2 U2373 ( .A(n2257), .B(n2280), .Z(n2258) );
  CND2X4 U2374 ( .A(n2259), .B(n2258), .Z(n2313) );
  CND2X4 U2375 ( .A(n2325), .B(n2345), .Z(n2386) );
  COND1X1 U2376 ( .A(n2389), .B(n2375), .C(n978), .Z(n2397) );
  COND1X1 U2377 ( .A(n2262), .B(n2373), .C(n2331), .Z(\req_vec_rr_d[10][2] )
         );
  CND2X4 U2378 ( .A(n2264), .B(n2263), .Z(n2384) );
  CND2X4 U2379 ( .A(n2266), .B(n2265), .Z(n2396) );
  COND1XL U2380 ( .A(n2379), .B(n2268), .C(n2267), .Z(n2269) );
  CNR2X1 U2381 ( .A(n2270), .B(n2269), .Z(n2275) );
  CND2X1 U2382 ( .A(n2271), .B(\req_vec_rr[11][3] ), .Z(n2272) );
  CND2IXL U2383 ( .B(n2277), .A(n2276), .Z(n2278) );
  CND3X1 U2384 ( .A(n977), .B(n2279), .C(n2278), .Z(n2281) );
  COR2X1 U2385 ( .A(n2348), .B(n2282), .Z(n2290) );
  CND2X1 U2386 ( .A(n2283), .B(\req_vec_rr[5][3] ), .Z(n2289) );
  CNR2XL U2387 ( .A(n2285), .B(n2284), .Z(n2288) );
  COND2X1 U2388 ( .A(n2352), .B(n2292), .C(n2371), .D(n2291), .Z(n2294) );
  CND3X2 U2389 ( .A(n2298), .B(n2297), .C(n2296), .Z(n2385) );
  CIVX2 U2390 ( .A(n2326), .Z(n2349) );
  CENX1 U2391 ( .A(n2361), .B(n2327), .Z(n2395) );
  COND1XL U2392 ( .A(n2299), .B(n2396), .C(n2395), .Z(\req_vec_rr_d[0][3] ) );
  CIVX4 U2393 ( .A(rst), .Z(n2412) );
  CNIVX4 U2394 ( .A(n2324), .Z(n2356) );
  COND1X1 U2395 ( .A(n2300), .B(n2356), .C(n2369), .Z(\req_vec_rr_d[12][0] )
         );
  COND1X1 U2396 ( .A(n2301), .B(n2373), .C(n2369), .Z(\req_vec_rr_d[2][0] ) );
  CNR2IX2 U2397 ( .B(n2326), .A(n2345), .Z(n2302) );
  CNR2X4 U2398 ( .A(n2389), .B(n2302), .Z(n2365) );
  CNIVX1 U2399 ( .A(n2416), .Z(n2308) );
  CIVDX3 U2400 ( .A(n2313), .Z0(n2325), .Z1(n2304) );
  CENX2 U2401 ( .A(n2358), .B(n2385), .Z(n2305) );
  CENX2 U2402 ( .A(n2305), .B(n2306), .Z(n2307) );
  CND2X2 U2403 ( .A(n2384), .B(n2307), .Z(n2309) );
  COND1X1 U2404 ( .A(n2308), .B(n2384), .C(n2309), .Z(\req_vec_rr_d[10][3] )
         );
  CIVX2 U2405 ( .A(n2309), .Z(n2311) );
  CNR2X2 U2406 ( .A(n2311), .B(n2310), .Z(n2417) );
  CNIVX1 U2407 ( .A(n2325), .Z(n2388) );
  CND2IX1 U2408 ( .B(n2396), .A(\req_vec_rr[11][2] ), .Z(n2312) );
  COAN1X1 U2409 ( .A(n918), .B(n2398), .C(n2369), .Z(n2420) );
  COAN1X1 U2410 ( .A(n922), .B(n2396), .C(n2369), .Z(n2419) );
  COAN1X1 U2411 ( .A(n920), .B(n2398), .C(n2369), .Z(n2421) );
  COAN1X1 U2412 ( .A(\req_vec_rr[11][3] ), .B(n2396), .C(n2347), .Z(
        \req_vec_rr_d[11][3] ) );
  COAN1X1 U2413 ( .A(n921), .B(n2396), .C(n2369), .Z(n2418) );
  CNIVX4 U2414 ( .A(n2324), .Z(n2373) );
  CIVX2 U2415 ( .A(n2314), .Z(n2315) );
  COND1X1 U2416 ( .A(n2315), .B(n2356), .C(n2369), .Z(\req_vec_rr_d[8][0] ) );
  COND1XL U2417 ( .A(n2317), .B(n2396), .C(n2388), .Z(\req_vec_rr_d[15][2] )
         );
  COAN1X1 U2418 ( .A(\req_vec_rr[7][2] ), .B(n2398), .C(n2318), .Z(n2406) );
  CENX2 U2419 ( .A(n2361), .B(n2386), .Z(n2387) );
  CIVX2 U2420 ( .A(n2387), .Z(n2383) );
  COND1X1 U2421 ( .A(n2323), .B(n2382), .C(n2369), .Z(\req_vec_rr_d[0][0] ) );
  CNIVX4 U2422 ( .A(n2324), .Z(n2382) );
  COND1X1 U2423 ( .A(n2328), .B(n2382), .C(n2370), .Z(\req_vec_rr_d[8][2] ) );
  COND1X1 U2424 ( .A(n2329), .B(n2382), .C(n2370), .Z(\req_vec_rr_d[0][2] ) );
  COND1X1 U2425 ( .A(n2330), .B(n2373), .C(n2365), .Z(\req_vec_rr_d[4][1] ) );
  COND1X1 U2426 ( .A(n2332), .B(n2373), .C(n2331), .Z(\req_vec_rr_d[2][2] ) );
  COND1X1 U2427 ( .A(n2333), .B(n2373), .C(n2365), .Z(\req_vec_rr_d[0][1] ) );
  COND1X1 U2428 ( .A(n2334), .B(n2356), .C(n2369), .Z(\req_vec_rr_d[6][0] ) );
  COND1X1 U2429 ( .A(n2335), .B(n2382), .C(n2365), .Z(\req_vec_rr_d[8][1] ) );
  COND1X1 U2430 ( .A(n2336), .B(n2382), .C(n2365), .Z(\req_vec_rr_d[12][1] )
         );
  COND1X1 U2431 ( .A(n2337), .B(n2382), .C(n917), .Z(\req_vec_rr_d[15][1] ) );
  CIVX2 U2432 ( .A(n2375), .Z(n2355) );
  CND2X1 U2433 ( .A(n2345), .B(n2340), .Z(n2341) );
  CAN2X1 U2434 ( .A(n2380), .B(n2341), .Z(n2409) );
  CND2X1 U2435 ( .A(n2345), .B(n2342), .Z(n2343) );
  CAN2X1 U2436 ( .A(n2380), .B(n2343), .Z(n2411) );
  CND2X1 U2437 ( .A(n2345), .B(n2344), .Z(n2346) );
  CAN2X1 U2438 ( .A(n2380), .B(n2346), .Z(n2410) );
  COND1X1 U2439 ( .A(n2348), .B(n2356), .C(n2347), .Z(\req_vec_rr_d[3][3] ) );
  CNR2X2 U2440 ( .A(n2349), .B(n2386), .Z(n2350) );
  CENX1 U2441 ( .A(n2361), .B(n2350), .Z(n2351) );
  COND1X1 U2442 ( .A(n2352), .B(n2373), .C(n2351), .Z(\req_vec_rr_d[6][3] ) );
  CENX1 U2443 ( .A(n2361), .B(n2353), .Z(n2368) );
  COND1X1 U2444 ( .A(n2354), .B(n2382), .C(n2368), .Z(\req_vec_rr_d[4][3] ) );
  COND1X1 U2445 ( .A(n2357), .B(n2373), .C(n2355), .Z(\req_vec_rr_d[9][2] ) );
  CENX1 U2446 ( .A(n2361), .B(n2358), .Z(n2378) );
  CIVX2 U2447 ( .A(n2378), .Z(n2359) );
  COND1X1 U2448 ( .A(n2360), .B(n2373), .C(n2359), .Z(\req_vec_rr_d[1][3] ) );
  CIVX1 U2449 ( .A(\req_vec_rr[15][3] ), .Z(n2362) );
  COND1X1 U2450 ( .A(n2362), .B(n2356), .C(n2361), .Z(\req_vec_rr_d[15][3] )
         );
  CND2X1 U2451 ( .A(n2365), .B(\req_vec_rr[10][1] ), .Z(n2363) );
  CND2X1 U2452 ( .A(n2367), .B(n2363), .Z(\req_vec_rr_d[10][1] ) );
  CND2X1 U2453 ( .A(n2365), .B(\req_vec_rr[14][1] ), .Z(n2364) );
  CND2X1 U2454 ( .A(n2367), .B(n2364), .Z(\req_vec_rr_d[14][1] ) );
  CND2X1 U2455 ( .A(n2365), .B(n926), .Z(n2366) );
  CND2X1 U2456 ( .A(n2367), .B(n2366), .Z(\req_vec_rr_d[6][1] ) );
  COAN1X1 U2457 ( .A(\req_vec_rr[11][0] ), .B(n2398), .C(n2369), .Z(n2407) );
  COAN1X1 U2458 ( .A(\req_vec_rr[12][2] ), .B(n2398), .C(n2370), .Z(
        \req_vec_rr_d[12][2] ) );
  COAN1X1 U2459 ( .A(\req_vec_rr[12][3] ), .B(n2396), .C(n2368), .Z(
        \req_vec_rr_d[12][3] ) );
  COAN1X1 U2460 ( .A(n919), .B(n2398), .C(n2369), .Z(n2408) );
  COAN1X1 U2461 ( .A(\req_vec_rr[4][2] ), .B(n2396), .C(n2370), .Z(
        \req_vec_rr_d[4][2] ) );
  COND1X1 U2462 ( .A(n2372), .B(n2382), .C(n2380), .Z(\req_vec_rr_d[5][1] ) );
  COND1X1 U2463 ( .A(n2374), .B(n2373), .C(n2380), .Z(\req_vec_rr_d[1][1] ) );
  CMXI2X1 U2464 ( .A0(n2376), .A1(n2394), .S(n2396), .Z(\req_vec_rr_d[13][2] )
         );
  CIVX2 U2465 ( .A(\req_vec_rr[13][3] ), .Z(n2377) );
  CMXI2X1 U2466 ( .A0(n2377), .A1(n2387), .S(n2396), .Z(\req_vec_rr_d[13][3] )
         );
  COND1X1 U2467 ( .A(n2381), .B(n2356), .C(n2380), .Z(\req_vec_rr_d[9][1] ) );
  CND2XL U2468 ( .A(n2386), .B(n2385), .Z(n2391) );
  CND3XL U2469 ( .A(n2389), .B(n2388), .C(n2387), .Z(n2390) );
  CND4X1 U2470 ( .A(n2393), .B(n2392), .C(n2391), .D(n2390), .Z(
        \req_vec_rr_d[14][3] ) );
  COAN1X1 U2471 ( .A(n923), .B(n2396), .C(n2395), .Z(\req_vec_rr_d[8][3] ) );
  CIVDX1 U2472 ( .A(n2397), .Z0(n2399), .Z1(n2331) );
  CMXI2X1 U2473 ( .A0(n1072), .A1(n2399), .S(n2398), .Z(\req_vec_rr_d[14][2] )
         );
  CMXI2X1 U2474 ( .A0(n2400), .A1(n2399), .S(n2398), .Z(\req_vec_rr_d[6][2] )
         );
endmodule

